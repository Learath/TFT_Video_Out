----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Sun Oct 26 17:57:07 2014
-- Parameters for CoreConfigMaster
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant DATA_LOCATION : integer := 256000;
end coreparameters;
