-- Version: v11.4 11.4.0.112

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_O2F                        : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC;

architecture DEF_ARCH of Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ_FAB
    port( A      : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_RCOSC_25_50MHZ_CLKINT, 
        \FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC <= 
        \FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\;

    I_RCOSC_25_50MHZ_FAB : RCOSC_25_50MHZ_FAB
      port map(A => 
        \FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\, 
        CLKOUT => N_RCOSC_25_50MHZ_CLKINT);
    
    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => 
        \FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    I_RCOSC_25_50MHZ_FAB_CLKINT : CLKINT
      port map(A => N_RCOSC_25_50MHZ_CLKINT, Y => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( HPMS_READY                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F                      : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0          : in    std_logic;
          INIT_DONE                                        : out   std_logic;
          POWER_ON_RESET_N                                 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : in    std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : in    std_logic;
          CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET     : in    std_logic;
          CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N         : out   std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \HPMS_READY\, 
        \sm0_areset_n_clk_base\, sm0_areset_n_clk_base_0, 
        \sm0_areset_n_rcosc\, sm0_areset_n_rcosc_0, 
        \count_ddr[0]_net_1\, \count_ddr_s[0]\, \ddr_settled\, 
        VCC_net_1, \un13_count_ddr\, GND_net_1, 
        \count_ddr_enable\, next_count_ddr_enable_0_sqmuxa, 
        \un1_next_ddr_ready_0_sqmuxa\, \mss_ready_select\, 
        \POWER_ON_RESET_N_clk_base\, N_6_i_0, 
        \sm0_state[0]_net_1\, \FDDR_CORE_RESET_N_int\, 
        \sm0_state[5]_net_1\, \mss_ready_state\, 
        \RESET_N_M2F_clk_base\, \sm0_state[6]_net_1\, 
        \sm0_state[4]_net_1\, \sm0_state_ns[2]_net_1\, 
        \sm0_state[3]_net_1\, \sm0_state_ns[3]_net_1\, 
        \sm0_state[2]_net_1\, \sm0_state_ns[4]_net_1\, 
        \sm0_state[1]_net_1\, \sm0_state_ns[5]_net_1\, 
        \sm0_state_ns_a3[6]_net_1\, sm0_areset_n_i_0_i, 
        sm0_areset_n_rcosc_q1, N_30_i_0, release_sdif3_core_q1, 
        release_sdif3_core, \POWER_ON_RESET_N_q1\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_q1\, 
        \sdif3_spll_lock_q1\, \count_ddr_enable_rcosc\, 
        \count_ddr_enable_q1\, \ddr_settled_clk_base\, 
        \ddr_settled_q1\, release_sdif3_core_clk_base, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \sm0_areset_n_q1\, 
        \CONFIG1_DONE_clk_base\, \CONFIG1_DONE_q1\, 
        \CONFIG2_DONE_clk_base\, \CONFIG2_DONE_q1\, 
        \sdif3_spll_lock_q2\, \count_ddr[1]_net_1\, 
        \count_ddr_s[1]\, \count_ddr[2]_net_1\, \count_ddr_s[2]\, 
        \count_ddr[3]_net_1\, \count_ddr_s[3]\, 
        \count_ddr[4]_net_1\, \count_ddr_s[4]\, 
        \count_ddr[5]_net_1\, \count_ddr_s[5]\, 
        \count_ddr[6]_net_1\, \count_ddr_s[6]\, 
        \count_ddr[7]_net_1\, \count_ddr_s[7]\, 
        \count_ddr[8]_net_1\, \count_ddr_s[8]_net_1\, 
        \count_ddr[9]_net_1\, \count_ddr_s[9]\, 
        \count_ddr[10]_net_1\, \count_ddr_s[10]\, 
        \count_ddr[11]_net_1\, \count_ddr_s[11]\, 
        \count_ddr[12]_net_1\, \count_ddr_s[12]\, 
        \count_ddr[13]_net_1\, \count_ddr_s[13]_net_1\, 
        \count_ddr_cry_1_FCO[12]\, \count_ddr_cry_3_FCO[12]\, 
        \count_ddr_cry[9]_net_1\, \count_ddr_cry[10]_net_1\, 
        \count_ddr_cry[11]_net_1\, \count_ddr_cry[12]_net_1\, 
        count_ddr_s_171_FCO, \count_ddr_cry[1]_net_1\, 
        \count_ddr_cry[2]_net_1\, \count_ddr_cry[3]_net_1\, 
        \count_ddr_cry[4]_net_1\, \count_ddr_cry[5]_net_1\, 
        \count_ddr_cry[6]_net_1\, \count_ddr_cry[7]_net_1\, 
        \un13_count_ddr_6\, \un8_ddr_settled_clk_base\, 
        \un13_count_ddr_9\, \un13_count_ddr_8\, 
        \un13_count_ddr_7\ : std_logic;

begin 

    HPMS_READY <= \HPMS_READY\;

    \sm0_state_ns[4]\ : CFG4
      generic map(INIT => x"FF70")

      port map(A => release_sdif3_core_clk_base, B => 
        \ddr_settled_clk_base\, C => \sm0_state[2]_net_1\, D => 
        next_count_ddr_enable_0_sqmuxa, Y => 
        \sm0_state_ns[4]_net_1\);
    
    sm0_areset_n_rcosc : SLE
      port map(D => sm0_areset_n_rcosc_q1, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_0_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_areset_n_rcosc\);
    
    \count_ddr[3]\ : SLE
      port map(D => \count_ddr_s[3]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[3]_net_1\);
    
    sm0_areset_n_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_i_0_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_areset_n_q1\);
    
    un13_count_ddr_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[7]_net_1\, B => 
        \count_ddr[6]_net_1\, C => \count_ddr[5]_net_1\, D => 
        \count_ddr[3]_net_1\, Y => \un13_count_ddr_8\);
    
    count_ddr_enable_q1 : SLE
      port map(D => \count_ddr_enable\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_rcosc_0, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_q1\);
    
    \sm0_state[6]\ : SLE
      port map(D => GND_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[6]_net_1\);
    
    count_ddr_s_171 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => count_ddr_s_171_FCO);
    
    sm0_areset_n_clk_base_RNIE6L5 : CLKINT
      port map(A => \sm0_areset_n_clk_base\, Y => 
        sm0_areset_n_clk_base_0);
    
    \sm0_state[2]\ : SLE
      port map(D => \sm0_state_ns[4]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[2]_net_1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    \count_ddr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[3]_net_1\, S => \count_ddr_s[4]\, Y => 
        OPEN, FCO => \count_ddr_cry[4]_net_1\);
    
    un8_ddr_settled_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \ddr_settled_clk_base\, B => 
        release_sdif3_core_clk_base, Y => 
        \un8_ddr_settled_clk_base\);
    
    INIT_DONE_int : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \sm0_state[0]_net_1\, ALn => sm0_areset_n_clk_base_0, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => INIT_DONE);
    
    \count_ddr[9]\ : SLE
      port map(D => \count_ddr_s[9]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[9]_net_1\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => N_30_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    
    count_ddr_enable_rcosc : SLE
      port map(D => \count_ddr_enable_q1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_rcosc_0, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_rcosc\);
    
    \count_ddr_cry_1[12]\ : ARI1
      generic map(INIT => x"48000")

      port map(A => \count_ddr[4]_net_1\, B => 
        \count_ddr[1]_net_1\, C => \count_ddr[2]_net_1\, D => 
        \count_ddr[3]_net_1\, FCI => \count_ddr[0]_net_1\, S => 
        OPEN, Y => OPEN, FCO => \count_ddr_cry_1_FCO[12]\);
    
    \count_ddr[7]\ : SLE
      port map(D => \count_ddr_s[7]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[7]_net_1\);
    
    \sm0_state_ns_a3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, Y => \sm0_state_ns_a3[6]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sm0_state[4]\ : SLE
      port map(D => \sm0_state_ns[2]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[4]_net_1\);
    
    MSS_HPMS_READY_int_RNO : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => N_30_i_0);
    
    un13_count_ddr_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \count_ddr[10]_net_1\, B => 
        \count_ddr[9]_net_1\, C => \count_ddr[8]_net_1\, D => 
        \count_ddr[4]_net_1\, Y => \un13_count_ddr_7\);
    
    count_ddr_enable : SLE
      port map(D => next_count_ddr_enable_0_sqmuxa, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_next_ddr_ready_0_sqmuxa\, ALn => 
        sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable\);
    
    \count_ddr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[9]_net_1\, S => \count_ddr_s[10]\, Y => 
        OPEN, FCO => \count_ddr_cry[10]_net_1\);
    
    \sm0_state[5]\ : SLE
      port map(D => \sm0_state[6]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[5]_net_1\);
    
    \count_ddr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[10]_net_1\, S => \count_ddr_s[11]\, Y => 
        OPEN, FCO => \count_ddr_cry[11]_net_1\);
    
    \count_ddr[8]\ : SLE
      port map(D => \count_ddr_s[8]_net_1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[8]_net_1\);
    
    \sm0_state_ns[2]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \CONFIG1_DONE_clk_base\, B => 
        \sm0_state[5]_net_1\, C => \sm0_state[4]_net_1\, Y => 
        \sm0_state_ns[2]_net_1\);
    
    sm0_areset_n_clk_base : SLE
      port map(D => \sm0_areset_n_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_i_0_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_areset_n_clk_base\);
    
    sm0_areset_n_rcosc_RNIK6M4 : CLKINT
      port map(A => \sm0_areset_n_rcosc\, Y => 
        sm0_areset_n_rcosc_0);
    
    \count_ddr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[11]_net_1\, S => \count_ddr_s[12]\, Y => 
        OPEN, FCO => \count_ddr_cry[12]_net_1\);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \sm0_state[1]\ : SLE
      port map(D => \sm0_state_ns[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[1]_net_1\);
    
    next_count_ddr_enable_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, Y => next_count_ddr_enable_0_sqmuxa);
    
    un13_count_ddr_6 : CFG2
      generic map(INIT => x"4")

      port map(A => \count_ddr[0]_net_1\, B => 
        \count_ddr[13]_net_1\, Y => \un13_count_ddr_6\);
    
    ddr_settled_clk_base : SLE
      port map(D => \ddr_settled_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_clk_base\);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FIC_2_APB_M_PRESET_N_q1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count_ddr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \count_ddr[0]_net_1\, Y => \count_ddr_s[0]\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => POWER_ON_RESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_clk_base\);
    
    \count_ddr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => count_ddr_s_171_FCO, S
         => \count_ddr_s[1]\, Y => OPEN, FCO => 
        \count_ddr_cry[1]_net_1\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_q1\);
    
    release_sdif0_core_q1 : SLE
      port map(D => release_sdif3_core, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        release_sdif3_core_q1);
    
    \count_ddr[10]\ : SLE
      port map(D => \count_ddr_s[10]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[10]_net_1\);
    
    \count_ddr_s[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[7]_net_1\, S => \count_ddr_s[8]_net_1\, Y
         => OPEN, FCO => OPEN);
    
    \count_ddr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[5]_net_1\, S => \count_ddr_s[6]\, Y => 
        OPEN, FCO => \count_ddr_cry[6]_net_1\);
    
    un13_count_ddr : CFG4
      generic map(INIT => x"8000")

      port map(A => \un13_count_ddr_8\, B => \un13_count_ddr_7\, 
        C => \un13_count_ddr_6\, D => \un13_count_ddr_9\, Y => 
        \un13_count_ddr\);
    
    MSS_HPMS_READY_int_RNIN6JD : CFG2
      generic map(INIT => x"8")

      port map(A => \HPMS_READY\, B => POWER_ON_RESET_N, Y => 
        sm0_areset_n_i_0_i);
    
    \count_ddr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[12]_net_1\, S => \count_ddr_s[13]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \count_ddr[5]\ : SLE
      port map(D => \count_ddr_s[5]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[5]_net_1\);
    
    \count_ddr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[2]_net_1\, S => \count_ddr_s[3]\, Y => 
        OPEN, FCO => \count_ddr_cry[3]_net_1\);
    
    \count_ddr[2]\ : SLE
      port map(D => \count_ddr_s[2]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[2]_net_1\);
    
    MSS_HPMS_READY_int_RNI3D17 : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => \HPMS_READY\);
    
    MDDR_DDR_AXI_S_CORE_RESET_N_0_a4 : CFG2
      generic map(INIT => x"4")

      port map(A => CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET, 
        B => \FDDR_CORE_RESET_N_int\, Y => 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N);
    
    sdif0_areset_n_rcosc_q1 : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_0_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => sm0_areset_n_rcosc_q1);
    
    \count_ddr[1]\ : SLE
      port map(D => \count_ddr_s[1]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[1]_net_1\);
    
    \sm0_state[0]\ : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \sm0_state_ns_a3[6]_net_1\, ALn => 
        sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[0]_net_1\);
    
    mss_ready_select_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => N_6_i_0);
    
    \count_ddr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[1]_net_1\, S => \count_ddr_s[2]\, Y => 
        OPEN, FCO => \count_ddr_cry[2]_net_1\);
    
    \count_ddr_cry_3[12]\ : ARI1
      generic map(INIT => x"48000")

      port map(A => \count_ddr[8]_net_1\, B => 
        \count_ddr[5]_net_1\, C => \count_ddr[6]_net_1\, D => 
        \count_ddr[7]_net_1\, FCI => \count_ddr_cry_1_FCO[12]\, S
         => OPEN, Y => OPEN, FCO => \count_ddr_cry_3_FCO[12]\);
    
    \count_ddr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[4]_net_1\, S => \count_ddr_s[5]\, Y => 
        OPEN, FCO => \count_ddr_cry[5]_net_1\);
    
    ddr_settled_q1 : SLE
      port map(D => \ddr_settled\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_q1\);
    
    \count_ddr[11]\ : SLE
      port map(D => \count_ddr_s[11]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[11]_net_1\);
    
    \sm0_state[3]\ : SLE
      port map(D => \sm0_state_ns[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[3]_net_1\);
    
    \sm0_state_ns[3]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \sm0_state[3]_net_1\, B => 
        \sdif3_spll_lock_q2\, C => \sm0_state[4]_net_1\, D => 
        \CONFIG1_DONE_clk_base\, Y => \sm0_state_ns[3]_net_1\);
    
    \count_ddr[0]\ : SLE
      port map(D => \count_ddr_s[0]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[0]_net_1\);
    
    CONFIG2_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG2_DONE, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_q1\);
    
    CONFIG2_DONE_clk_base : SLE
      port map(D => \CONFIG2_DONE_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_clk_base\);
    
    CONFIG1_DONE_clk_base : SLE
      port map(D => \CONFIG1_DONE_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_6_i_0, 
        ALn => \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \count_ddr[4]\ : SLE
      port map(D => \count_ddr_s[4]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[4]_net_1\);
    
    \count_ddr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[6]_net_1\, S => \count_ddr_s[7]\, Y => 
        OPEN, FCO => \count_ddr_cry[7]_net_1\);
    
    un13_count_ddr_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[12]_net_1\, B => 
        \count_ddr[11]_net_1\, C => \count_ddr[2]_net_1\, D => 
        \count_ddr[1]_net_1\, Y => \un13_count_ddr_9\);
    
    release_sdif0_core : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => sm0_areset_n_rcosc_0, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => release_sdif3_core);
    
    FDDR_CORE_RESET_N_int : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \sm0_state[5]_net_1\, ALn => sm0_areset_n_clk_base_0, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FDDR_CORE_RESET_N_int\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => POWER_ON_RESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_q1\);
    
    \count_ddr[12]\ : SLE
      port map(D => \count_ddr_s[12]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[12]_net_1\);
    
    ddr_settled : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => \un13_count_ddr\, ALn => sm0_areset_n_rcosc_0, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ddr_settled\);
    
    \count_ddr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry_3_FCO[12]\, S => \count_ddr_s[9]\, Y => 
        OPEN, FCO => \count_ddr_cry[9]_net_1\);
    
    \count_ddr[6]\ : SLE
      port map(D => \count_ddr_s[6]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[6]_net_1\);
    
    CONFIG1_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG1_DONE, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_q1\);
    
    sdif3_spll_lock_q1 : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sdif3_spll_lock_q1\);
    
    release_sdif0_core_clk_base : SLE
      port map(D => release_sdif3_core_q1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        release_sdif3_core_clk_base);
    
    sdif3_spll_lock_q2 : SLE
      port map(D => \sdif3_spll_lock_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => sm0_areset_n_clk_base_0, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sdif3_spll_lock_q2\);
    
    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    un1_next_ddr_ready_0_sqmuxa : CFG4
      generic map(INIT => x"F888")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, C => \ddr_settled_clk_base\, D => 
        \sm0_state[2]_net_1\, Y => \un1_next_ddr_ready_0_sqmuxa\);
    
    \count_ddr[13]\ : SLE
      port map(D => \count_ddr_s[13]_net_1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => sm0_areset_n_rcosc_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[13]_net_1\);
    
    \sm0_state_ns[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, C => \un8_ddr_settled_clk_base\, D
         => \sm0_state[2]_net_1\, Y => \sm0_state_ns[5]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Igloo2_TFT_Video_Out_Test_HPMS is

    port( MDDR_DQS                                                    : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                                     : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DM_RDQS                                                : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_BA                                                     : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                                   : out   std_logic_vector(15 downto 0);
          xhdl1328_i_m_0_1                                            : in    std_logic_vector(0 to 0);
          ConfigMaster_0_M_HRDATA                                     : out   std_logic_vector(31 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA                         : out   std_logic_vector(15 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR                             : in    std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE                             : in    std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HTRANS                            : in    std_logic_vector(1 to 1);
          CoreAHBLite_1_AHBmslave16_HWDATA                            : in    std_logic_vector(31 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR                          : in    std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA                         : in    std_logic_vector(15 downto 0);
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_0  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_1  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_2  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_3  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_4  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_5  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_6  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_7  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_8  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_9  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_10 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_11 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_12 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_13 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_14 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_15 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_16 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18 : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                                : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                                    : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i_0                                : out   std_logic;
          MDDR_WE_N                                                   : out   std_logic;
          MDDR_RESET_N                                                : out   std_logic;
          MDDR_RAS_N                                                  : out   std_logic;
          MDDR_ODT                                                    : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                                       : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                                        : in    std_logic;
          MDDR_CS_N                                                   : out   std_logic;
          MDDR_CKE                                                    : out   std_logic;
          MDDR_CAS_N                                                  : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY                            : inout std_logic := 'Z';
          CoreAHBLite_1_AHBmslave16_HREADY_i_m                        : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F            : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx     : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE    : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY                         : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR                        : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx                             : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE                            : in    std_logic;
          HPMS_DDR_FIC_SUBSYSTEM_LOCK                                 : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY    : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR   : in    std_logic;
          CORECONFIGP_0_SOFT_RESET_F2M_i_0                            : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0                     : in    std_logic;
          CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N                    : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE                        : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx                          : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE                         : in    std_logic;
          MDDR_CLK_N                                                  : out   std_logic;
          MDDR_CLK                                                    : out   std_logic
        );

end Igloo2_TFT_Video_Out_Test_HPMS;

architecture DEF_ARCH of Igloo2_TFT_Video_Out_Test_HPMS is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MSS_010

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := "");

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OUTBUF_DIFF
    generic (IOSTD:string := "");

    port( D    : in    std_logic := 'U';
          PADP : out   std_logic;
          PADN : out   std_logic
        );
  end component;

    signal CONFIG_PRESET_N, \CORECONFIGP_0_APB_S_PRESET_N\, 
        FIC_2_APB_M_PCLK, \CORECONFIGP_0_APB_S_PCLK\, 
        MSS_ADLIB_INST_DRAM_WEN, MSS_ADLIB_INST_DRAM_RSTN, 
        MSS_ADLIB_INST_DRAM_RASN, MSS_ADLIB_INST_DRAM_ODT, 
        \DRAM_FIFO_WE_OUT_net_0[0]\, MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        MDDR_DQS_1_PAD_Y, \DRAM_DQS_OUT_net_0[1]\, 
        \DRAM_DQS_OE_net_0[1]\, MDDR_DQS_0_PAD_Y, 
        \DRAM_DQS_OUT_net_0[0]\, \DRAM_DQS_OE_net_0[0]\, 
        MDDR_DQ_15_PAD_Y, \DRAM_DQ_OUT_net_0[15]\, 
        \DRAM_DQ_OE_net_0[15]\, MDDR_DQ_14_PAD_Y, 
        \DRAM_DQ_OUT_net_0[14]\, \DRAM_DQ_OE_net_0[14]\, 
        MDDR_DQ_13_PAD_Y, \DRAM_DQ_OUT_net_0[13]\, 
        \DRAM_DQ_OE_net_0[13]\, MDDR_DQ_12_PAD_Y, 
        \DRAM_DQ_OUT_net_0[12]\, \DRAM_DQ_OE_net_0[12]\, 
        MDDR_DQ_11_PAD_Y, \DRAM_DQ_OUT_net_0[11]\, 
        \DRAM_DQ_OE_net_0[11]\, MDDR_DQ_10_PAD_Y, 
        \DRAM_DQ_OUT_net_0[10]\, \DRAM_DQ_OE_net_0[10]\, 
        MDDR_DQ_9_PAD_Y, \DRAM_DQ_OUT_net_0[9]\, 
        \DRAM_DQ_OE_net_0[9]\, MDDR_DQ_8_PAD_Y, 
        \DRAM_DQ_OUT_net_0[8]\, \DRAM_DQ_OE_net_0[8]\, 
        MDDR_DQ_7_PAD_Y, \DRAM_DQ_OUT_net_0[7]\, 
        \DRAM_DQ_OE_net_0[7]\, MDDR_DQ_6_PAD_Y, 
        \DRAM_DQ_OUT_net_0[6]\, \DRAM_DQ_OE_net_0[6]\, 
        MDDR_DQ_5_PAD_Y, \DRAM_DQ_OUT_net_0[5]\, 
        \DRAM_DQ_OE_net_0[5]\, MDDR_DQ_4_PAD_Y, 
        \DRAM_DQ_OUT_net_0[4]\, \DRAM_DQ_OE_net_0[4]\, 
        MDDR_DQ_3_PAD_Y, \DRAM_DQ_OUT_net_0[3]\, 
        \DRAM_DQ_OE_net_0[3]\, MDDR_DQ_2_PAD_Y, 
        \DRAM_DQ_OUT_net_0[2]\, \DRAM_DQ_OE_net_0[2]\, 
        MDDR_DQ_1_PAD_Y, \DRAM_DQ_OUT_net_0[1]\, 
        \DRAM_DQ_OE_net_0[1]\, MDDR_DQ_0_PAD_Y, 
        \DRAM_DQ_OUT_net_0[0]\, \DRAM_DQ_OE_net_0[0]\, 
        MDDR_DM_RDQS_1_PAD_Y, \DRAM_DM_RDQS_OUT_net_0[1]\, 
        \DM_OE_net_0[1]\, MDDR_DM_RDQS_0_PAD_Y, 
        \DRAM_DM_RDQS_OUT_net_0[0]\, \DM_OE_net_0[0]\, 
        MSS_ADLIB_INST_DRAM_CSN, MSS_ADLIB_INST_DRAM_CKE, 
        MSS_ADLIB_INST_DRAM_CASN, \DRAM_BA_net_0[2]\, 
        \DRAM_BA_net_0[1]\, \DRAM_BA_net_0[0]\, 
        \DRAM_ADDR_net_0[15]\, \DRAM_ADDR_net_0[14]\, 
        \DRAM_ADDR_net_0[13]\, \DRAM_ADDR_net_0[12]\, 
        \DRAM_ADDR_net_0[11]\, \DRAM_ADDR_net_0[10]\, 
        \DRAM_ADDR_net_0[9]\, \DRAM_ADDR_net_0[8]\, 
        \DRAM_ADDR_net_0[7]\, \DRAM_ADDR_net_0[6]\, 
        \DRAM_ADDR_net_0[5]\, \DRAM_ADDR_net_0[4]\, 
        \DRAM_ADDR_net_0[3]\, \DRAM_ADDR_net_0[2]\, 
        \DRAM_ADDR_net_0[1]\, \DRAM_ADDR_net_0[0]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[0]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[1]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[2]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[3]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[4]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[5]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[6]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[7]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[8]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[9]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[10]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[11]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[12]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[13]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[14]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[15]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[16]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[17]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[18]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[19]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[20]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[21]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[22]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[25]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[26]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[28]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[30]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[31]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[24]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[27]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[29]\, 
        \CoreAHBLite_1_AHBmslave16_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave0_HREADY, VCC_net_1, GND_net_1, 
        MSS_ADLIB_INST_DRAM_CLK : std_logic;
    signal nc228, nc203, nc216, nc194, nc151, nc23, nc175, nc58, 
        nc116, nc74, nc133, nc238, nc167, nc84, nc39, nc72, nc212, 
        nc205, nc82, nc145, nc181, nc160, nc57, nc156, nc125, 
        nc211, nc73, nc107, nc66, nc83, nc9, nc171, nc54, nc135, 
        nc41, nc100, nc52, nc186, nc29, nc118, nc60, nc141, nc193, 
        nc214, nc45, nc53, nc121, nc176, nc220, nc158, nc209, 
        nc162, nc11, nc131, nc96, nc79, nc226, nc146, nc230, nc89, 
        nc119, nc48, nc213, nc126, nc195, nc188, nc15, nc236, 
        nc102, nc3, nc207, nc47, nc90, nc222, nc159, nc136, nc178, 
        nc215, nc59, nc221, nc232, nc18, nc44, nc117, nc189, 
        nc164, nc148, nc42, nc231, nc191, nc17, nc2, nc110, nc128, 
        nc43, nc179, nc157, nc36, nc224, nc61, nc104, nc138, nc14, 
        nc150, nc196, nc234, nc149, nc12, nc219, nc30, nc187, 
        nc65, nc7, nc129, nc8, nc223, nc13, nc180, nc26, nc177, 
        nc139, nc233, nc163, nc112, nc68, nc49, nc217, nc170, 
        nc91, nc225, nc5, nc20, nc198, nc147, nc67, nc152, nc127, 
        nc103, nc235, nc76, nc208, nc140, nc86, nc95, nc120, 
        nc165, nc137, nc64, nc19, nc70, nc182, nc62, nc199, nc80, 
        nc130, nc98, nc114, nc56, nc105, nc63, nc172, nc229, nc97, 
        nc161, nc31, nc154, nc50, nc142, nc94, nc197, nc122, nc35, 
        nc4, nc227, nc92, nc101, nc184, nc200, nc190, nc166, 
        nc132, nc21, nc237, nc93, nc69, nc206, nc174, nc38, nc113, 
        nc218, nc106, nc25, nc1, nc37, nc202, nc144, nc153, nc46, 
        nc71, nc124, nc81, nc201, nc168, nc34, nc28, nc115, nc192, 
        nc134, nc32, nc40, nc99, nc75, nc183, nc85, nc27, nc108, 
        nc16, nc155, nc51, nc33, nc204, nc173, nc169, nc78, nc24, 
        nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, nc77, 
        nc6, nc109, nc87, nc123 : std_logic;

begin 

    CORECONFIGP_0_APB_S_PRESET_N <= 
        \CORECONFIGP_0_APB_S_PRESET_N\;
    CORECONFIGP_0_APB_S_PCLK <= \CORECONFIGP_0_APB_S_PCLK\;

    MDDR_ADDR_6_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[6]\, PAD => MDDR_ADDR(6));
    
    MSS_ADLIB_INST_RNIHJLG_9 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[10]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(10));
    
    MDDR_CAS_N_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CASN, PAD => MDDR_CAS_N);
    
    MSS_ADLIB_INST_RNIHJLG_2 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[3]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(3));
    
    MDDR_RESET_N_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_RSTN, PAD => MDDR_RESET_N);
    
    MDDR_ODT_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_ODT, PAD => MDDR_ODT);
    
    MSS_ADLIB_INST_RNIHJLG_29 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[30]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(30));
    
    MDDR_ADDR_11_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[11]\, PAD => MDDR_ADDR(11));
    
    MSS_ADLIB_INST_RNIHJLG_11 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[12]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(12));
    
    MDDR_DQ_10_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(10), D => \DRAM_DQ_OUT_net_0[10]\, 
        E => \DRAM_DQ_OE_net_0[10]\, Y => MDDR_DQ_10_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_7 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[8]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(8));
    
    MSS_ADLIB_INST_RNIHJLG_31 : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        xhdl1328_i_m_0_1(0), Y => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m);
    
    MDDR_DQ_1_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(1), D => \DRAM_DQ_OUT_net_0[1]\, E
         => \DRAM_DQ_OE_net_0[1]\, Y => MDDR_DQ_1_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_16 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[17]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(17));
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIU0V1_0 : CFG1
      generic map(INIT => "01")

      port map(A => \CORECONFIGP_0_APB_S_PCLK\, Y => 
        CORECONFIGP_0_APB_S_PCLK_i_0);
    
    MSS_ADLIB_INST_RNIHJLG_13 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[14]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(14));
    
    MDDR_ADDR_7_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[7]\, PAD => MDDR_ADDR(7));
    
    MDDR_DQ_11_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(11), D => \DRAM_DQ_OUT_net_0[11]\, 
        E => \DRAM_DQ_OE_net_0[11]\, Y => MDDR_DQ_11_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_21 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[22]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(22));
    
    MDDR_DQ_9_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(9), D => \DRAM_DQ_OUT_net_0[9]\, E
         => \DRAM_DQ_OE_net_0[9]\, Y => MDDR_DQ_9_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_26 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[27]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(27));
    
    MDDR_DQ_3_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(3), D => \DRAM_DQ_OUT_net_0[3]\, E
         => \DRAM_DQ_OE_net_0[3]\, Y => MDDR_DQ_3_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_23 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[24]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(24));
    
    MDDR_DQ_0_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(0), D => \DRAM_DQ_OUT_net_0[0]\, E
         => \DRAM_DQ_OE_net_0[0]\, Y => MDDR_DQ_0_PAD_Y);
    
    MDDR_ADDR_12_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[12]\, PAD => MDDR_ADDR(12));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MDDR_DQ_2_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(2), D => \DRAM_DQ_OUT_net_0[2]\, E
         => \DRAM_DQ_OE_net_0[2]\, Y => MDDR_DQ_2_PAD_Y);
    
    MDDR_DQ_12_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(12), D => \DRAM_DQ_OUT_net_0[12]\, 
        E => \DRAM_DQ_OE_net_0[12]\, Y => MDDR_DQ_12_PAD_Y);
    
    MDDR_CKE_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CKE, PAD => MDDR_CKE);
    
    MDDR_ADDR_2_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[2]\, PAD => MDDR_ADDR(2));
    
    MDDR_ADDR_13_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[13]\, PAD => MDDR_ADDR(13));
    
    MDDR_ADDR_5_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[5]\, PAD => MDDR_ADDR(5));
    
    MDDR_DM_RDQS_1_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DM_RDQS(1), D => 
        \DRAM_DM_RDQS_OUT_net_0[1]\, E => \DM_OE_net_0[1]\, Y => 
        MDDR_DM_RDQS_1_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_17 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[18]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(18));
    
    MDDR_DQS_0_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQS(0), D => \DRAM_DQS_OUT_net_0[0]\, 
        E => \DRAM_DQS_OE_net_0[0]\, Y => MDDR_DQS_0_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_14 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[15]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(15));
    
    MDDR_DQS_1_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQS(1), D => \DRAM_DQS_OUT_net_0[1]\, 
        E => \DRAM_DQS_OE_net_0[1]\, Y => MDDR_DQS_1_PAD_Y);
    
    MDDR_DQ_15_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(15), D => \DRAM_DQ_OUT_net_0[15]\, 
        E => \DRAM_DQ_OE_net_0[15]\, Y => MDDR_DQ_15_PAD_Y);
    
    MDDR_DM_RDQS_0_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DM_RDQS(0), D => 
        \DRAM_DM_RDQS_OUT_net_0[0]\, E => \DM_OE_net_0[0]\, Y => 
        MDDR_DM_RDQS_0_PAD_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNIHJLG_27 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[28]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(28));
    
    MSS_ADLIB_INST_RNIHJLG_24 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[25]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(25));
    
    MDDR_DQ_8_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(8), D => \DRAM_DQ_OUT_net_0[8]\, E
         => \DRAM_DQ_OE_net_0[8]\, Y => MDDR_DQ_8_PAD_Y);
    
    MDDR_ADDR_9_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[9]\, PAD => MDDR_ADDR(9));
    
    MDDR_BA_2_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_BA_net_0[2]\, PAD => MDDR_BA(2));
    
    MDDR_ADDR_14_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[14]\, PAD => MDDR_ADDR(14));
    
    MSS_ADLIB_INST_RNIHJLG_8 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[9]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(9));
    
    MSS_ADLIB_INST_RNIHJLG_5 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[6]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(6));
    
    MSS_ADLIB_INST : MSS_010

              generic map(INIT => "00" & x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C31D00820000608EC0000003FFFFE400000010000000000000000F11C0000007EDFFC010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem")

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => FIC_2_APB_M_PCLK, COMMS_INT
         => OPEN, CONFIG_PRESET_N => CONFIG_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc216, EDAC_ERROR(4) => nc194, 
        EDAC_ERROR(3) => nc151, EDAC_ERROR(2) => nc23, 
        EDAC_ERROR(1) => nc175, EDAC_ERROR(0) => nc58, 
        F_FM0_RDATA(31) => \CoreAHBLite_1_AHBmslave16_HRDATA[31]\, 
        F_FM0_RDATA(30) => \CoreAHBLite_1_AHBmslave16_HRDATA[30]\, 
        F_FM0_RDATA(29) => \CoreAHBLite_1_AHBmslave16_HRDATA[29]\, 
        F_FM0_RDATA(28) => \CoreAHBLite_1_AHBmslave16_HRDATA[28]\, 
        F_FM0_RDATA(27) => \CoreAHBLite_1_AHBmslave16_HRDATA[27]\, 
        F_FM0_RDATA(26) => \CoreAHBLite_1_AHBmslave16_HRDATA[26]\, 
        F_FM0_RDATA(25) => \CoreAHBLite_1_AHBmslave16_HRDATA[25]\, 
        F_FM0_RDATA(24) => \CoreAHBLite_1_AHBmslave16_HRDATA[24]\, 
        F_FM0_RDATA(23) => \CoreAHBLite_1_AHBmslave16_HRDATA[23]\, 
        F_FM0_RDATA(22) => \CoreAHBLite_1_AHBmslave16_HRDATA[22]\, 
        F_FM0_RDATA(21) => \CoreAHBLite_1_AHBmslave16_HRDATA[21]\, 
        F_FM0_RDATA(20) => \CoreAHBLite_1_AHBmslave16_HRDATA[20]\, 
        F_FM0_RDATA(19) => \CoreAHBLite_1_AHBmslave16_HRDATA[19]\, 
        F_FM0_RDATA(18) => \CoreAHBLite_1_AHBmslave16_HRDATA[18]\, 
        F_FM0_RDATA(17) => \CoreAHBLite_1_AHBmslave16_HRDATA[17]\, 
        F_FM0_RDATA(16) => \CoreAHBLite_1_AHBmslave16_HRDATA[16]\, 
        F_FM0_RDATA(15) => \CoreAHBLite_1_AHBmslave16_HRDATA[15]\, 
        F_FM0_RDATA(14) => \CoreAHBLite_1_AHBmslave16_HRDATA[14]\, 
        F_FM0_RDATA(13) => \CoreAHBLite_1_AHBmslave16_HRDATA[13]\, 
        F_FM0_RDATA(12) => \CoreAHBLite_1_AHBmslave16_HRDATA[12]\, 
        F_FM0_RDATA(11) => \CoreAHBLite_1_AHBmslave16_HRDATA[11]\, 
        F_FM0_RDATA(10) => \CoreAHBLite_1_AHBmslave16_HRDATA[10]\, 
        F_FM0_RDATA(9) => \CoreAHBLite_1_AHBmslave16_HRDATA[9]\, 
        F_FM0_RDATA(8) => \CoreAHBLite_1_AHBmslave16_HRDATA[8]\, 
        F_FM0_RDATA(7) => \CoreAHBLite_1_AHBmslave16_HRDATA[7]\, 
        F_FM0_RDATA(6) => \CoreAHBLite_1_AHBmslave16_HRDATA[6]\, 
        F_FM0_RDATA(5) => \CoreAHBLite_1_AHBmslave16_HRDATA[5]\, 
        F_FM0_RDATA(4) => \CoreAHBLite_1_AHBmslave16_HRDATA[4]\, 
        F_FM0_RDATA(3) => \CoreAHBLite_1_AHBmslave16_HRDATA[3]\, 
        F_FM0_RDATA(2) => \CoreAHBLite_1_AHBmslave16_HRDATA[2]\, 
        F_FM0_RDATA(1) => \CoreAHBLite_1_AHBmslave16_HRDATA[1]\, 
        F_FM0_RDATA(0) => \CoreAHBLite_1_AHBmslave16_HRDATA[0]\, 
        F_FM0_READYOUT => CoreAHBLite_1_AHBmslave16_HREADY, 
        F_FM0_RESP => OPEN, F_HM0_ADDR(31) => nc116, 
        F_HM0_ADDR(30) => nc74, F_HM0_ADDR(29) => nc133, 
        F_HM0_ADDR(28) => nc238, F_HM0_ADDR(27) => nc167, 
        F_HM0_ADDR(26) => nc84, F_HM0_ADDR(25) => nc39, 
        F_HM0_ADDR(24) => nc72, F_HM0_ADDR(23) => nc212, 
        F_HM0_ADDR(22) => nc205, F_HM0_ADDR(21) => nc82, 
        F_HM0_ADDR(20) => nc145, F_HM0_ADDR(19) => nc181, 
        F_HM0_ADDR(18) => nc160, F_HM0_ADDR(17) => nc57, 
        F_HM0_ADDR(16) => nc156, F_HM0_ADDR(15) => nc125, 
        F_HM0_ADDR(14) => nc211, F_HM0_ADDR(13) => nc73, 
        F_HM0_ADDR(12) => nc107, F_HM0_ADDR(11) => nc66, 
        F_HM0_ADDR(10) => nc83, F_HM0_ADDR(9) => nc9, 
        F_HM0_ADDR(8) => nc171, F_HM0_ADDR(7) => nc54, 
        F_HM0_ADDR(6) => nc135, F_HM0_ADDR(5) => nc41, 
        F_HM0_ADDR(4) => nc100, F_HM0_ADDR(3) => nc52, 
        F_HM0_ADDR(2) => nc186, F_HM0_ADDR(1) => nc29, 
        F_HM0_ADDR(0) => nc118, F_HM0_ENABLE => OPEN, F_HM0_SEL
         => OPEN, F_HM0_SIZE(1) => nc60, F_HM0_SIZE(0) => nc141, 
        F_HM0_TRANS1 => OPEN, F_HM0_WDATA(31) => nc193, 
        F_HM0_WDATA(30) => nc214, F_HM0_WDATA(29) => nc45, 
        F_HM0_WDATA(28) => nc53, F_HM0_WDATA(27) => nc121, 
        F_HM0_WDATA(26) => nc176, F_HM0_WDATA(25) => nc220, 
        F_HM0_WDATA(24) => nc158, F_HM0_WDATA(23) => nc209, 
        F_HM0_WDATA(22) => nc162, F_HM0_WDATA(21) => nc11, 
        F_HM0_WDATA(20) => nc131, F_HM0_WDATA(19) => nc96, 
        F_HM0_WDATA(18) => nc79, F_HM0_WDATA(17) => nc226, 
        F_HM0_WDATA(16) => nc146, F_HM0_WDATA(15) => nc230, 
        F_HM0_WDATA(14) => nc89, F_HM0_WDATA(13) => nc119, 
        F_HM0_WDATA(12) => nc48, F_HM0_WDATA(11) => nc213, 
        F_HM0_WDATA(10) => nc126, F_HM0_WDATA(9) => nc195, 
        F_HM0_WDATA(8) => nc188, F_HM0_WDATA(7) => nc15, 
        F_HM0_WDATA(6) => nc236, F_HM0_WDATA(5) => nc102, 
        F_HM0_WDATA(4) => nc3, F_HM0_WDATA(3) => nc207, 
        F_HM0_WDATA(2) => nc47, F_HM0_WDATA(1) => nc90, 
        F_HM0_WDATA(0) => nc222, F_HM0_WRITE => OPEN, 
        FAB_CHRGVBUS => OPEN, FAB_DISCHRGVBUS => OPEN, 
        FAB_DMPULLDOWN => OPEN, FAB_DPPULLDOWN => OPEN, 
        FAB_DRVVBUS => OPEN, FAB_IDPULLUP => OPEN, FAB_OPMODE(1)
         => nc159, FAB_OPMODE(0) => nc136, FAB_SUSPENDM => OPEN, 
        FAB_TERMSEL => OPEN, FAB_TXVALID => OPEN, FAB_VCONTROL(3)
         => nc178, FAB_VCONTROL(2) => nc215, FAB_VCONTROL(1) => 
        nc59, FAB_VCONTROL(0) => nc221, FAB_VCONTROLLOADM => OPEN, 
        FAB_XCVRSEL(1) => nc232, FAB_XCVRSEL(0) => nc18, 
        FAB_XDATAOUT(7) => nc44, FAB_XDATAOUT(6) => nc117, 
        FAB_XDATAOUT(5) => nc189, FAB_XDATAOUT(4) => nc164, 
        FAB_XDATAOUT(3) => nc148, FAB_XDATAOUT(2) => nc42, 
        FAB_XDATAOUT(1) => nc231, FAB_XDATAOUT(0) => nc191, 
        FACC_GLMUX_SEL => OPEN, FIC32_0_MASTER(1) => nc17, 
        FIC32_0_MASTER(0) => nc2, FIC32_1_MASTER(1) => nc110, 
        FIC32_1_MASTER(0) => nc128, FPGA_RESET_N => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, GTX_CLK
         => OPEN, H2F_INTERRUPT(15) => nc43, H2F_INTERRUPT(14)
         => nc179, H2F_INTERRUPT(13) => nc157, H2F_INTERRUPT(12)
         => nc36, H2F_INTERRUPT(11) => nc224, H2F_INTERRUPT(10)
         => nc61, H2F_INTERRUPT(9) => nc104, H2F_INTERRUPT(8) => 
        nc138, H2F_INTERRUPT(7) => nc14, H2F_INTERRUPT(6) => 
        nc150, H2F_INTERRUPT(5) => nc196, H2F_INTERRUPT(4) => 
        nc234, H2F_INTERRUPT(3) => nc149, H2F_INTERRUPT(2) => 
        nc12, H2F_INTERRUPT(1) => nc219, H2F_INTERRUPT(0) => nc30, 
        H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_A => OPEN, I2C1_SDA_MGPIO0A_H2F_B
         => OPEN, MDCF => OPEN, MDOENF => OPEN, MDOF => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13, 
        PER2_FABRIC_PADDR(14) => nc187, PER2_FABRIC_PADDR(13) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11, 
        PER2_FABRIC_PADDR(12) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10, 
        PER2_FABRIC_PADDR(11) => nc65, PER2_FABRIC_PADDR(10) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8, 
        PER2_FABRIC_PADDR(9) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7, 
        PER2_FABRIC_PADDR(8) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6, 
        PER2_FABRIC_PADDR(7) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5, 
        PER2_FABRIC_PADDR(6) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4, 
        PER2_FABRIC_PADDR(5) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3, 
        PER2_FABRIC_PADDR(4) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        PER2_FABRIC_PADDR(3) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        PER2_FABRIC_PADDR(2) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        PER2_FABRIC_PENABLE => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        PER2_FABRIC_PSEL => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx, 
        PER2_FABRIC_PWDATA(31) => nc7, PER2_FABRIC_PWDATA(30) => 
        nc129, PER2_FABRIC_PWDATA(29) => nc8, 
        PER2_FABRIC_PWDATA(28) => nc223, PER2_FABRIC_PWDATA(27)
         => nc13, PER2_FABRIC_PWDATA(26) => nc180, 
        PER2_FABRIC_PWDATA(25) => nc26, PER2_FABRIC_PWDATA(24)
         => nc177, PER2_FABRIC_PWDATA(23) => nc139, 
        PER2_FABRIC_PWDATA(22) => nc233, PER2_FABRIC_PWDATA(21)
         => nc163, PER2_FABRIC_PWDATA(20) => nc112, 
        PER2_FABRIC_PWDATA(19) => nc68, PER2_FABRIC_PWDATA(18)
         => nc49, PER2_FABRIC_PWDATA(17) => nc217, 
        PER2_FABRIC_PWDATA(16) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_16, 
        PER2_FABRIC_PWDATA(15) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_15, 
        PER2_FABRIC_PWDATA(14) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_14, 
        PER2_FABRIC_PWDATA(13) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_13, 
        PER2_FABRIC_PWDATA(12) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_12, 
        PER2_FABRIC_PWDATA(11) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_11, 
        PER2_FABRIC_PWDATA(10) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_10, 
        PER2_FABRIC_PWDATA(9) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_9, 
        PER2_FABRIC_PWDATA(8) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_8, 
        PER2_FABRIC_PWDATA(7) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_7, 
        PER2_FABRIC_PWDATA(6) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_6, 
        PER2_FABRIC_PWDATA(5) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_5, 
        PER2_FABRIC_PWDATA(4) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_4, 
        PER2_FABRIC_PWDATA(3) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_3, 
        PER2_FABRIC_PWDATA(2) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_2, 
        PER2_FABRIC_PWDATA(1) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_1, 
        PER2_FABRIC_PWDATA(0) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_0, 
        PER2_FABRIC_PWRITE => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        RTC_MATCH => OPEN, SLEEPDEEP => OPEN, SLEEPHOLDACK => 
        OPEN, SLEEPING => OPEN, SMBALERT_NO0 => OPEN, 
        SMBALERT_NO1 => OPEN, SMBSUS_NO0 => OPEN, SMBSUS_NO1 => 
        OPEN, SPI0_CLK_OUT => OPEN, SPI0_SDI_MGPIO5A_H2F_A => 
        OPEN, SPI0_SDI_MGPIO5A_H2F_B => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_A => OPEN, SPI0_SDO_MGPIO6A_H2F_B
         => OPEN, SPI0_SS0_MGPIO7A_H2F_A => OPEN, 
        SPI0_SS0_MGPIO7A_H2F_B => OPEN, SPI0_SS1_MGPIO8A_H2F_A
         => OPEN, SPI0_SS1_MGPIO8A_H2F_B => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_A => OPEN, SPI0_SS2_MGPIO9A_H2F_B
         => OPEN, SPI0_SS3_MGPIO10A_H2F_A => OPEN, 
        SPI0_SS3_MGPIO10A_H2F_B => OPEN, SPI0_SS4_MGPIO19A_H2F_A
         => OPEN, SPI0_SS5_MGPIO20A_H2F_A => OPEN, 
        SPI0_SS6_MGPIO21A_H2F_A => OPEN, SPI0_SS7_MGPIO22A_H2F_A
         => OPEN, SPI1_CLK_OUT => OPEN, SPI1_SDI_MGPIO11A_H2F_A
         => OPEN, SPI1_SDI_MGPIO11A_H2F_B => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_A => OPEN, SPI1_SDO_MGPIO12A_H2F_B
         => OPEN, SPI1_SS0_MGPIO13A_H2F_A => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_B => OPEN, SPI1_SS1_MGPIO14A_H2F_A
         => OPEN, SPI1_SS1_MGPIO14A_H2F_B => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_A => OPEN, SPI1_SS2_MGPIO15A_H2F_B
         => OPEN, SPI1_SS3_MGPIO16A_H2F_A => OPEN, 
        SPI1_SS3_MGPIO16A_H2F_B => OPEN, SPI1_SS4_MGPIO17A_H2F_A
         => OPEN, SPI1_SS5_MGPIO18A_H2F_A => OPEN, 
        SPI1_SS6_MGPIO23A_H2F_A => OPEN, SPI1_SS7_MGPIO24A_H2F_A
         => OPEN, TCGF(9) => nc170, TCGF(8) => nc91, TCGF(7) => 
        nc225, TCGF(6) => nc5, TCGF(5) => nc20, TCGF(4) => nc198, 
        TCGF(3) => nc147, TCGF(2) => nc67, TCGF(1) => nc152, 
        TCGF(0) => nc127, TRACECLK => OPEN, TRACEDATA(3) => nc103, 
        TRACEDATA(2) => nc235, TRACEDATA(1) => nc76, TRACEDATA(0)
         => nc208, TX_CLK => OPEN, TX_ENF => OPEN, TX_ERRF => 
        OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc140, 
        TXD_RIF(2) => nc86, TXD_RIF(1) => nc95, TXD_RIF(0) => 
        nc120, TXDF(7) => nc165, TXDF(6) => nc137, TXDF(5) => 
        nc64, TXDF(4) => nc19, TXDF(3) => nc70, TXDF(2) => nc182, 
        TXDF(1) => nc62, TXDF(0) => nc199, TXEV => OPEN, 
        WDOGTIMEOUT => OPEN, F_ARREADY_HREADYOUT1 => OPEN, 
        F_AWREADY_HREADYOUT0 => CoreAHBLite_0_AHBmslave0_HREADY, 
        F_BID(3) => nc80, F_BID(2) => nc130, F_BID(1) => nc98, 
        F_BID(0) => nc114, F_BRESP_HRESP0(1) => nc56, 
        F_BRESP_HRESP0(0) => nc105, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc63, F_RDATA_HRDATA01(62) => 
        nc172, F_RDATA_HRDATA01(61) => nc229, 
        F_RDATA_HRDATA01(60) => nc97, F_RDATA_HRDATA01(59) => 
        nc161, F_RDATA_HRDATA01(58) => nc31, F_RDATA_HRDATA01(57)
         => nc154, F_RDATA_HRDATA01(56) => nc50, 
        F_RDATA_HRDATA01(55) => nc142, F_RDATA_HRDATA01(54) => 
        nc94, F_RDATA_HRDATA01(53) => nc197, F_RDATA_HRDATA01(52)
         => nc122, F_RDATA_HRDATA01(51) => nc35, 
        F_RDATA_HRDATA01(50) => nc4, F_RDATA_HRDATA01(49) => 
        nc227, F_RDATA_HRDATA01(48) => nc92, F_RDATA_HRDATA01(47)
         => nc101, F_RDATA_HRDATA01(46) => nc184, 
        F_RDATA_HRDATA01(45) => nc200, F_RDATA_HRDATA01(44) => 
        nc190, F_RDATA_HRDATA01(43) => nc166, 
        F_RDATA_HRDATA01(42) => nc132, F_RDATA_HRDATA01(41) => 
        nc21, F_RDATA_HRDATA01(40) => nc237, F_RDATA_HRDATA01(39)
         => nc93, F_RDATA_HRDATA01(38) => nc69, 
        F_RDATA_HRDATA01(37) => nc206, F_RDATA_HRDATA01(36) => 
        nc174, F_RDATA_HRDATA01(35) => nc38, F_RDATA_HRDATA01(34)
         => nc113, F_RDATA_HRDATA01(33) => nc218, 
        F_RDATA_HRDATA01(32) => nc106, F_RDATA_HRDATA01(31) => 
        nc25, F_RDATA_HRDATA01(30) => nc1, F_RDATA_HRDATA01(29)
         => nc37, F_RDATA_HRDATA01(28) => nc202, 
        F_RDATA_HRDATA01(27) => nc144, F_RDATA_HRDATA01(26) => 
        nc153, F_RDATA_HRDATA01(25) => nc46, F_RDATA_HRDATA01(24)
         => nc71, F_RDATA_HRDATA01(23) => nc124, 
        F_RDATA_HRDATA01(22) => nc81, F_RDATA_HRDATA01(21) => 
        nc201, F_RDATA_HRDATA01(20) => nc168, 
        F_RDATA_HRDATA01(19) => nc34, F_RDATA_HRDATA01(18) => 
        nc28, F_RDATA_HRDATA01(17) => nc115, F_RDATA_HRDATA01(16)
         => nc192, F_RDATA_HRDATA01(15) => nc134, 
        F_RDATA_HRDATA01(14) => nc32, F_RDATA_HRDATA01(13) => 
        nc40, F_RDATA_HRDATA01(12) => nc99, F_RDATA_HRDATA01(11)
         => nc75, F_RDATA_HRDATA01(10) => nc183, 
        F_RDATA_HRDATA01(9) => nc85, F_RDATA_HRDATA01(8) => nc27, 
        F_RDATA_HRDATA01(7) => nc108, F_RDATA_HRDATA01(6) => nc16, 
        F_RDATA_HRDATA01(5) => nc155, F_RDATA_HRDATA01(4) => nc51, 
        F_RDATA_HRDATA01(3) => nc33, F_RDATA_HRDATA01(2) => nc204, 
        F_RDATA_HRDATA01(1) => nc173, F_RDATA_HRDATA01(0) => 
        nc169, F_RID(3) => nc78, F_RID(2) => nc24, F_RID(1) => 
        nc88, F_RID(0) => nc111, F_RLAST => OPEN, 
        F_RRESP_HRESP1(1) => nc55, F_RRESP_HRESP1(0) => nc10, 
        F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), 
        MDDR_FABRIC_PRDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), 
        MDDR_FABRIC_PRDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), 
        MDDR_FABRIC_PRDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), 
        MDDR_FABRIC_PRDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), 
        MDDR_FABRIC_PRDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), 
        MDDR_FABRIC_PRDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), 
        MDDR_FABRIC_PRDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), 
        MDDR_FABRIC_PRDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), 
        MDDR_FABRIC_PRDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), 
        MDDR_FABRIC_PRDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), 
        MDDR_FABRIC_PRDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), 
        MDDR_FABRIC_PRDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), 
        MDDR_FABRIC_PRDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), 
        MDDR_FABRIC_PRDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), 
        MDDR_FABRIC_PRDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), 
        MDDR_FABRIC_PREADY => CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        MDDR_FABRIC_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        CoreAHBLite_1_AHBmslave16_HADDR(31), F_FM0_ADDR(30) => 
        CoreAHBLite_1_AHBmslave16_HADDR(30), F_FM0_ADDR(29) => 
        CoreAHBLite_1_AHBmslave16_HADDR(29), F_FM0_ADDR(28) => 
        CoreAHBLite_1_AHBmslave16_HADDR(28), F_FM0_ADDR(27) => 
        CoreAHBLite_1_AHBmslave16_HADDR(27), F_FM0_ADDR(26) => 
        CoreAHBLite_1_AHBmslave16_HADDR(26), F_FM0_ADDR(25) => 
        CoreAHBLite_1_AHBmslave16_HADDR(25), F_FM0_ADDR(24) => 
        CoreAHBLite_1_AHBmslave16_HADDR(24), F_FM0_ADDR(23) => 
        CoreAHBLite_1_AHBmslave16_HADDR(23), F_FM0_ADDR(22) => 
        CoreAHBLite_1_AHBmslave16_HADDR(22), F_FM0_ADDR(21) => 
        CoreAHBLite_1_AHBmslave16_HADDR(21), F_FM0_ADDR(20) => 
        CoreAHBLite_1_AHBmslave16_HADDR(20), F_FM0_ADDR(19) => 
        CoreAHBLite_1_AHBmslave16_HADDR(19), F_FM0_ADDR(18) => 
        CoreAHBLite_1_AHBmslave16_HADDR(18), F_FM0_ADDR(17) => 
        CoreAHBLite_1_AHBmslave16_HADDR(17), F_FM0_ADDR(16) => 
        CoreAHBLite_1_AHBmslave16_HADDR(16), F_FM0_ADDR(15) => 
        CoreAHBLite_1_AHBmslave16_HADDR(15), F_FM0_ADDR(14) => 
        CoreAHBLite_1_AHBmslave16_HADDR(14), F_FM0_ADDR(13) => 
        CoreAHBLite_1_AHBmslave16_HADDR(13), F_FM0_ADDR(12) => 
        CoreAHBLite_1_AHBmslave16_HADDR(12), F_FM0_ADDR(11) => 
        CoreAHBLite_1_AHBmslave16_HADDR(11), F_FM0_ADDR(10) => 
        CoreAHBLite_1_AHBmslave16_HADDR(10), F_FM0_ADDR(9) => 
        CoreAHBLite_1_AHBmslave16_HADDR(9), F_FM0_ADDR(8) => 
        CoreAHBLite_1_AHBmslave16_HADDR(8), F_FM0_ADDR(7) => 
        CoreAHBLite_1_AHBmslave16_HADDR(7), F_FM0_ADDR(6) => 
        CoreAHBLite_1_AHBmslave16_HADDR(6), F_FM0_ADDR(5) => 
        CoreAHBLite_1_AHBmslave16_HADDR(5), F_FM0_ADDR(4) => 
        CoreAHBLite_1_AHBmslave16_HADDR(4), F_FM0_ADDR(3) => 
        CoreAHBLite_1_AHBmslave16_HADDR(3), F_FM0_ADDR(2) => 
        CoreAHBLite_1_AHBmslave16_HADDR(2), F_FM0_ADDR(1) => 
        CoreAHBLite_1_AHBmslave16_HADDR(1), F_FM0_ADDR(0) => 
        CoreAHBLite_1_AHBmslave16_HADDR(0), F_FM0_ENABLE => 
        GND_net_1, F_FM0_MASTLOCK => GND_net_1, F_FM0_READY => 
        CoreAHBLite_1_AHBmslave16_HREADY, F_FM0_SEL => 
        CoreAHBLite_1_AHBmslave16_HSELx, F_FM0_SIZE(1) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(1), F_FM0_SIZE(0) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(0), F_FM0_TRANS1 => 
        CoreAHBLite_1_AHBmslave16_HTRANS(1), F_FM0_WDATA(31) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(31), F_FM0_WDATA(30) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(30), F_FM0_WDATA(29) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(29), F_FM0_WDATA(28) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(28), F_FM0_WDATA(27) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(27), F_FM0_WDATA(26) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(26), F_FM0_WDATA(25) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(25), F_FM0_WDATA(24) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(24), F_FM0_WDATA(23) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(23), F_FM0_WDATA(22) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(22), F_FM0_WDATA(21) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(21), F_FM0_WDATA(20) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(20), F_FM0_WDATA(19) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(19), F_FM0_WDATA(18) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(18), F_FM0_WDATA(17) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(17), F_FM0_WDATA(16) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(16), F_FM0_WDATA(15) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(15), F_FM0_WDATA(14) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(14), F_FM0_WDATA(13) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(13), F_FM0_WDATA(12) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(12), F_FM0_WDATA(11) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(11), F_FM0_WDATA(10) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(10), F_FM0_WDATA(9) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(9), F_FM0_WDATA(8) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(8), F_FM0_WDATA(7) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(7), F_FM0_WDATA(6) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(6), F_FM0_WDATA(5) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(5), F_FM0_WDATA(4) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(4), F_FM0_WDATA(3) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(3), F_FM0_WDATA(2) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(2), F_FM0_WDATA(1) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(1), F_FM0_WDATA(0) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(0), F_FM0_WRITE => 
        CoreAHBLite_1_AHBmslave16_HWRITE, F_HM0_RDATA(31) => 
        GND_net_1, F_HM0_RDATA(30) => GND_net_1, F_HM0_RDATA(29)
         => GND_net_1, F_HM0_RDATA(28) => GND_net_1, 
        F_HM0_RDATA(27) => GND_net_1, F_HM0_RDATA(26) => 
        GND_net_1, F_HM0_RDATA(25) => GND_net_1, F_HM0_RDATA(24)
         => GND_net_1, F_HM0_RDATA(23) => GND_net_1, 
        F_HM0_RDATA(22) => GND_net_1, F_HM0_RDATA(21) => 
        GND_net_1, F_HM0_RDATA(20) => GND_net_1, F_HM0_RDATA(19)
         => GND_net_1, F_HM0_RDATA(18) => GND_net_1, 
        F_HM0_RDATA(17) => GND_net_1, F_HM0_RDATA(16) => 
        GND_net_1, F_HM0_RDATA(15) => GND_net_1, F_HM0_RDATA(14)
         => GND_net_1, F_HM0_RDATA(13) => GND_net_1, 
        F_HM0_RDATA(12) => GND_net_1, F_HM0_RDATA(11) => 
        GND_net_1, F_HM0_RDATA(10) => GND_net_1, F_HM0_RDATA(9)
         => GND_net_1, F_HM0_RDATA(8) => GND_net_1, 
        F_HM0_RDATA(7) => GND_net_1, F_HM0_RDATA(6) => GND_net_1, 
        F_HM0_RDATA(5) => GND_net_1, F_HM0_RDATA(4) => GND_net_1, 
        F_HM0_RDATA(3) => GND_net_1, F_HM0_RDATA(2) => GND_net_1, 
        F_HM0_RDATA(1) => GND_net_1, F_HM0_RDATA(0) => GND_net_1, 
        F_HM0_READY => VCC_net_1, F_HM0_RESP => GND_net_1, 
        FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, 
        FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        GND_net_1, FAB_PLL_LOCK => HPMS_DDR_FIC_SUBSYSTEM_LOCK, 
        FAB_RXACTIVE => VCC_net_1, FAB_RXERROR => VCC_net_1, 
        FAB_RXVALID => VCC_net_1, FAB_RXVALIDH => GND_net_1, 
        FAB_SESSEND => VCC_net_1, FAB_TXREADY => VCC_net_1, 
        FAB_VBUSVALID => VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, 
        FAB_VSTATUS(6) => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => VCC_net_1, 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => VCC_net_1, 
        MGPIO30B_F2H_GPIN => VCC_net_1, MGPIO31B_F2H_GPIN => 
        VCC_net_1, MGPIO3A_F2H_GPIN => VCC_net_1, 
        MGPIO4A_F2H_GPIN => VCC_net_1, MGPIO5A_F2H_GPIN => 
        VCC_net_1, MGPIO6A_F2H_GPIN => VCC_net_1, 
        MGPIO7A_F2H_GPIN => VCC_net_1, MGPIO8A_F2H_GPIN => 
        VCC_net_1, MGPIO9A_F2H_GPIN => VCC_net_1, 
        MMUART0_CTS_F2H_SCP => VCC_net_1, MMUART0_DCD_F2H_SCP => 
        VCC_net_1, MMUART0_DSR_F2H_SCP => VCC_net_1, 
        MMUART0_DTR_F2H_SCP => VCC_net_1, MMUART0_RI_F2H_SCP => 
        VCC_net_1, MMUART0_RTS_F2H_SCP => VCC_net_1, 
        MMUART0_RXD_F2H_SCP => VCC_net_1, MMUART0_SCK_F2H_SCP => 
        VCC_net_1, MMUART0_TXD_F2H_SCP => VCC_net_1, 
        MMUART1_CTS_F2H_SCP => VCC_net_1, MMUART1_DCD_F2H_SCP => 
        VCC_net_1, MMUART1_DSR_F2H_SCP => VCC_net_1, 
        MMUART1_RI_F2H_SCP => VCC_net_1, MMUART1_RTS_F2H_SCP => 
        VCC_net_1, MMUART1_RXD_F2H_SCP => VCC_net_1, 
        MMUART1_SCK_F2H_SCP => VCC_net_1, MMUART1_TXD_F2H_SCP => 
        VCC_net_1, PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18, 
        PER2_FABRIC_PRDATA(17) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18, 
        PER2_FABRIC_PRDATA(16) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16, 
        PER2_FABRIC_PRDATA(15) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15, 
        PER2_FABRIC_PRDATA(14) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14, 
        PER2_FABRIC_PRDATA(13) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13, 
        PER2_FABRIC_PRDATA(12) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12, 
        PER2_FABRIC_PRDATA(11) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11, 
        PER2_FABRIC_PRDATA(10) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10, 
        PER2_FABRIC_PRDATA(9) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9, 
        PER2_FABRIC_PRDATA(8) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8, 
        PER2_FABRIC_PRDATA(7) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7, 
        PER2_FABRIC_PRDATA(6) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6, 
        PER2_FABRIC_PRDATA(5) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5, 
        PER2_FABRIC_PRDATA(4) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4, 
        PER2_FABRIC_PRDATA(3) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3, 
        PER2_FABRIC_PRDATA(2) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2, 
        PER2_FABRIC_PRDATA(1) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1, 
        PER2_FABRIC_PRDATA(0) => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0, 
        PER2_FABRIC_PREADY => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY, 
        PER2_FABRIC_PSLVERR => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR, 
        RCGF(9) => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => 
        VCC_net_1, RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, 
        RCGF(4) => VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => 
        VCC_net_1, RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, 
        RX_CLKPF => VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => 
        VCC_net_1, RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, 
        RXDF(6) => VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => 
        VCC_net_1, RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, 
        RXDF(1) => VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ
         => GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1
         => VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => CORECONFIGP_0_SOFT_RESET_F2M_i_0, 
        XCLK_FAB => VCC_net_1, CLK_BASE => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, CLK_MDDR_APB => 
        \CORECONFIGP_0_APB_S_PCLK\, F_ARADDR_HADDR1(31) => 
        VCC_net_1, F_ARADDR_HADDR1(30) => VCC_net_1, 
        F_ARADDR_HADDR1(29) => VCC_net_1, F_ARADDR_HADDR1(28) => 
        VCC_net_1, F_ARADDR_HADDR1(27) => VCC_net_1, 
        F_ARADDR_HADDR1(26) => VCC_net_1, F_ARADDR_HADDR1(25) => 
        VCC_net_1, F_ARADDR_HADDR1(24) => VCC_net_1, 
        F_ARADDR_HADDR1(23) => VCC_net_1, F_ARADDR_HADDR1(22) => 
        VCC_net_1, F_ARADDR_HADDR1(21) => VCC_net_1, 
        F_ARADDR_HADDR1(20) => VCC_net_1, F_ARADDR_HADDR1(19) => 
        VCC_net_1, F_ARADDR_HADDR1(18) => VCC_net_1, 
        F_ARADDR_HADDR1(17) => VCC_net_1, F_ARADDR_HADDR1(16) => 
        VCC_net_1, F_ARADDR_HADDR1(15) => VCC_net_1, 
        F_ARADDR_HADDR1(14) => VCC_net_1, F_ARADDR_HADDR1(13) => 
        VCC_net_1, F_ARADDR_HADDR1(12) => VCC_net_1, 
        F_ARADDR_HADDR1(11) => VCC_net_1, F_ARADDR_HADDR1(10) => 
        VCC_net_1, F_ARADDR_HADDR1(9) => VCC_net_1, 
        F_ARADDR_HADDR1(8) => VCC_net_1, F_ARADDR_HADDR1(7) => 
        VCC_net_1, F_ARADDR_HADDR1(6) => VCC_net_1, 
        F_ARADDR_HADDR1(5) => VCC_net_1, F_ARADDR_HADDR1(4) => 
        VCC_net_1, F_ARADDR_HADDR1(3) => VCC_net_1, 
        F_ARADDR_HADDR1(2) => VCC_net_1, F_ARADDR_HADDR1(1) => 
        VCC_net_1, F_ARADDR_HADDR1(0) => VCC_net_1, 
        F_ARBURST_HTRANS1(1) => GND_net_1, F_ARBURST_HTRANS1(0)
         => GND_net_1, F_ARID_HSEL1(3) => GND_net_1, 
        F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1) => 
        GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => GND_net_1, F_AWADDR_HADDR0(30) => 
        GND_net_1, F_AWADDR_HADDR0(29) => GND_net_1, 
        F_AWADDR_HADDR0(28) => GND_net_1, F_AWADDR_HADDR0(27) => 
        GND_net_1, F_AWADDR_HADDR0(26) => GND_net_1, 
        F_AWADDR_HADDR0(25) => GND_net_1, F_AWADDR_HADDR0(24) => 
        GND_net_1, F_AWADDR_HADDR0(23) => GND_net_1, 
        F_AWADDR_HADDR0(22) => GND_net_1, F_AWADDR_HADDR0(21) => 
        GND_net_1, F_AWADDR_HADDR0(20) => GND_net_1, 
        F_AWADDR_HADDR0(19) => GND_net_1, F_AWADDR_HADDR0(18) => 
        GND_net_1, F_AWADDR_HADDR0(17) => GND_net_1, 
        F_AWADDR_HADDR0(16) => GND_net_1, F_AWADDR_HADDR0(15) => 
        GND_net_1, F_AWADDR_HADDR0(14) => GND_net_1, 
        F_AWADDR_HADDR0(13) => GND_net_1, F_AWADDR_HADDR0(12) => 
        GND_net_1, F_AWADDR_HADDR0(11) => GND_net_1, 
        F_AWADDR_HADDR0(10) => GND_net_1, F_AWADDR_HADDR0(9) => 
        GND_net_1, F_AWADDR_HADDR0(8) => GND_net_1, 
        F_AWADDR_HADDR0(7) => GND_net_1, F_AWADDR_HADDR0(6) => 
        GND_net_1, F_AWADDR_HADDR0(5) => GND_net_1, 
        F_AWADDR_HADDR0(4) => GND_net_1, F_AWADDR_HADDR0(3) => 
        GND_net_1, F_AWADDR_HADDR0(2) => GND_net_1, 
        F_AWADDR_HADDR0(1) => GND_net_1, F_AWADDR_HADDR0(0) => 
        GND_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => GND_net_1, 
        F_WDATA_HWDATA01(30) => GND_net_1, F_WDATA_HWDATA01(29)
         => GND_net_1, F_WDATA_HWDATA01(28) => GND_net_1, 
        F_WDATA_HWDATA01(27) => GND_net_1, F_WDATA_HWDATA01(26)
         => GND_net_1, F_WDATA_HWDATA01(25) => GND_net_1, 
        F_WDATA_HWDATA01(24) => GND_net_1, F_WDATA_HWDATA01(23)
         => GND_net_1, F_WDATA_HWDATA01(22) => GND_net_1, 
        F_WDATA_HWDATA01(21) => GND_net_1, F_WDATA_HWDATA01(20)
         => GND_net_1, F_WDATA_HWDATA01(19) => GND_net_1, 
        F_WDATA_HWDATA01(18) => GND_net_1, F_WDATA_HWDATA01(17)
         => GND_net_1, F_WDATA_HWDATA01(16) => GND_net_1, 
        F_WDATA_HWDATA01(15) => GND_net_1, F_WDATA_HWDATA01(14)
         => GND_net_1, F_WDATA_HWDATA01(13) => GND_net_1, 
        F_WDATA_HWDATA01(12) => GND_net_1, F_WDATA_HWDATA01(11)
         => GND_net_1, F_WDATA_HWDATA01(10) => GND_net_1, 
        F_WDATA_HWDATA01(9) => GND_net_1, F_WDATA_HWDATA01(8) => 
        GND_net_1, F_WDATA_HWDATA01(7) => GND_net_1, 
        F_WDATA_HWDATA01(6) => GND_net_1, F_WDATA_HWDATA01(5) => 
        GND_net_1, F_WDATA_HWDATA01(4) => GND_net_1, 
        F_WDATA_HWDATA01(3) => GND_net_1, F_WDATA_HWDATA01(2) => 
        GND_net_1, F_WDATA_HWDATA01(1) => GND_net_1, 
        F_WDATA_HWDATA01(0) => GND_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        CoreAHBLite_0_AHBmslave0_HREADY, F_WLAST => GND_net_1, 
        F_WSTRB(7) => GND_net_1, F_WSTRB(6) => GND_net_1, 
        F_WSTRB(5) => GND_net_1, F_WSTRB(4) => GND_net_1, 
        F_WSTRB(3) => GND_net_1, F_WSTRB(2) => GND_net_1, 
        F_WSTRB(1) => GND_net_1, F_WSTRB(0) => GND_net_1, 
        F_WVALID => GND_net_1, FPGA_MDDR_ARESET_N => 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N, 
        MDDR_FABRIC_PADDR(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10), 
        MDDR_FABRIC_PADDR(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9), 
        MDDR_FABRIC_PADDR(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8), 
        MDDR_FABRIC_PADDR(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7), 
        MDDR_FABRIC_PADDR(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6), 
        MDDR_FABRIC_PADDR(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5), 
        MDDR_FABRIC_PADDR(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4), 
        MDDR_FABRIC_PADDR(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3), 
        MDDR_FABRIC_PADDR(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2), 
        MDDR_FABRIC_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, MDDR_FABRIC_PSEL
         => CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        MDDR_FABRIC_PWDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15), 
        MDDR_FABRIC_PWDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14), 
        MDDR_FABRIC_PWDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13), 
        MDDR_FABRIC_PWDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12), 
        MDDR_FABRIC_PWDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11), 
        MDDR_FABRIC_PWDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10), 
        MDDR_FABRIC_PWDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9), 
        MDDR_FABRIC_PWDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8), 
        MDDR_FABRIC_PWDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7), 
        MDDR_FABRIC_PWDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6), 
        MDDR_FABRIC_PWDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5), 
        MDDR_FABRIC_PWDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4), 
        MDDR_FABRIC_PWDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3), 
        MDDR_FABRIC_PWDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2), 
        MDDR_FABRIC_PWDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1), 
        MDDR_FABRIC_PWDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0), 
        MDDR_FABRIC_PWRITE => CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        PRESET_N => \CORECONFIGP_0_APB_S_PRESET_N\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => MDDR_DM_RDQS_1_PAD_Y, DM_IN(0)
         => MDDR_DM_RDQS_0_PAD_Y, DRAM_DQ_IN(17) => GND_net_1, 
        DRAM_DQ_IN(16) => GND_net_1, DRAM_DQ_IN(15) => 
        MDDR_DQ_15_PAD_Y, DRAM_DQ_IN(14) => MDDR_DQ_14_PAD_Y, 
        DRAM_DQ_IN(13) => MDDR_DQ_13_PAD_Y, DRAM_DQ_IN(12) => 
        MDDR_DQ_12_PAD_Y, DRAM_DQ_IN(11) => MDDR_DQ_11_PAD_Y, 
        DRAM_DQ_IN(10) => MDDR_DQ_10_PAD_Y, DRAM_DQ_IN(9) => 
        MDDR_DQ_9_PAD_Y, DRAM_DQ_IN(8) => MDDR_DQ_8_PAD_Y, 
        DRAM_DQ_IN(7) => MDDR_DQ_7_PAD_Y, DRAM_DQ_IN(6) => 
        MDDR_DQ_6_PAD_Y, DRAM_DQ_IN(5) => MDDR_DQ_5_PAD_Y, 
        DRAM_DQ_IN(4) => MDDR_DQ_4_PAD_Y, DRAM_DQ_IN(3) => 
        MDDR_DQ_3_PAD_Y, DRAM_DQ_IN(2) => MDDR_DQ_2_PAD_Y, 
        DRAM_DQ_IN(1) => MDDR_DQ_1_PAD_Y, DRAM_DQ_IN(0) => 
        MDDR_DQ_0_PAD_Y, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => MDDR_DQS_1_PAD_Y, DRAM_DQS_IN(0) => 
        MDDR_DQS_0_PAD_Y, DRAM_FIFO_WE_IN(1) => GND_net_1, 
        DRAM_FIFO_WE_IN(0) => MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => GND_net_1, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => GND_net_1, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => GND_net_1, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => GND_net_1, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, SPI1_SCK_IN
         => GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => \DRAM_ADDR_net_0[15]\, DRAM_ADDR(14) => 
        \DRAM_ADDR_net_0[14]\, DRAM_ADDR(13) => 
        \DRAM_ADDR_net_0[13]\, DRAM_ADDR(12) => 
        \DRAM_ADDR_net_0[12]\, DRAM_ADDR(11) => 
        \DRAM_ADDR_net_0[11]\, DRAM_ADDR(10) => 
        \DRAM_ADDR_net_0[10]\, DRAM_ADDR(9) => 
        \DRAM_ADDR_net_0[9]\, DRAM_ADDR(8) => 
        \DRAM_ADDR_net_0[8]\, DRAM_ADDR(7) => 
        \DRAM_ADDR_net_0[7]\, DRAM_ADDR(6) => 
        \DRAM_ADDR_net_0[6]\, DRAM_ADDR(5) => 
        \DRAM_ADDR_net_0[5]\, DRAM_ADDR(4) => 
        \DRAM_ADDR_net_0[4]\, DRAM_ADDR(3) => 
        \DRAM_ADDR_net_0[3]\, DRAM_ADDR(2) => 
        \DRAM_ADDR_net_0[2]\, DRAM_ADDR(1) => 
        \DRAM_ADDR_net_0[1]\, DRAM_ADDR(0) => 
        \DRAM_ADDR_net_0[0]\, DRAM_BA(2) => \DRAM_BA_net_0[2]\, 
        DRAM_BA(1) => \DRAM_BA_net_0[1]\, DRAM_BA(0) => 
        \DRAM_BA_net_0[0]\, DRAM_CASN => MSS_ADLIB_INST_DRAM_CASN, 
        DRAM_CKE => MSS_ADLIB_INST_DRAM_CKE, DRAM_CLK => 
        MSS_ADLIB_INST_DRAM_CLK, DRAM_CSN => 
        MSS_ADLIB_INST_DRAM_CSN, DRAM_DM_RDQS_OUT(2) => nc22, 
        DRAM_DM_RDQS_OUT(1) => \DRAM_DM_RDQS_OUT_net_0[1]\, 
        DRAM_DM_RDQS_OUT(0) => \DRAM_DM_RDQS_OUT_net_0[0]\, 
        DRAM_DQ_OUT(17) => nc210, DRAM_DQ_OUT(16) => nc185, 
        DRAM_DQ_OUT(15) => \DRAM_DQ_OUT_net_0[15]\, 
        DRAM_DQ_OUT(14) => \DRAM_DQ_OUT_net_0[14]\, 
        DRAM_DQ_OUT(13) => \DRAM_DQ_OUT_net_0[13]\, 
        DRAM_DQ_OUT(12) => \DRAM_DQ_OUT_net_0[12]\, 
        DRAM_DQ_OUT(11) => \DRAM_DQ_OUT_net_0[11]\, 
        DRAM_DQ_OUT(10) => \DRAM_DQ_OUT_net_0[10]\, 
        DRAM_DQ_OUT(9) => \DRAM_DQ_OUT_net_0[9]\, DRAM_DQ_OUT(8)
         => \DRAM_DQ_OUT_net_0[8]\, DRAM_DQ_OUT(7) => 
        \DRAM_DQ_OUT_net_0[7]\, DRAM_DQ_OUT(6) => 
        \DRAM_DQ_OUT_net_0[6]\, DRAM_DQ_OUT(5) => 
        \DRAM_DQ_OUT_net_0[5]\, DRAM_DQ_OUT(4) => 
        \DRAM_DQ_OUT_net_0[4]\, DRAM_DQ_OUT(3) => 
        \DRAM_DQ_OUT_net_0[3]\, DRAM_DQ_OUT(2) => 
        \DRAM_DQ_OUT_net_0[2]\, DRAM_DQ_OUT(1) => 
        \DRAM_DQ_OUT_net_0[1]\, DRAM_DQ_OUT(0) => 
        \DRAM_DQ_OUT_net_0[0]\, DRAM_DQS_OUT(2) => nc143, 
        DRAM_DQS_OUT(1) => \DRAM_DQS_OUT_net_0[1]\, 
        DRAM_DQS_OUT(0) => \DRAM_DQS_OUT_net_0[0]\, 
        DRAM_FIFO_WE_OUT(1) => nc77, DRAM_FIFO_WE_OUT(0) => 
        \DRAM_FIFO_WE_OUT_net_0[0]\, DRAM_ODT => 
        MSS_ADLIB_INST_DRAM_ODT, DRAM_RASN => 
        MSS_ADLIB_INST_DRAM_RASN, DRAM_RSTN => 
        MSS_ADLIB_INST_DRAM_RSTN, DRAM_WEN => 
        MSS_ADLIB_INST_DRAM_WEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, SPI1_SCK_OUT
         => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => OPEN, 
        SPI1_SS5_MGPIO18A_OUT => OPEN, SPI1_SS6_MGPIO23A_OUT => 
        OPEN, SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => 
        OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc6, 
        DM_OE(1) => \DM_OE_net_0[1]\, DM_OE(0) => 
        \DM_OE_net_0[0]\, DRAM_DQ_OE(17) => nc109, DRAM_DQ_OE(16)
         => nc87, DRAM_DQ_OE(15) => \DRAM_DQ_OE_net_0[15]\, 
        DRAM_DQ_OE(14) => \DRAM_DQ_OE_net_0[14]\, DRAM_DQ_OE(13)
         => \DRAM_DQ_OE_net_0[13]\, DRAM_DQ_OE(12) => 
        \DRAM_DQ_OE_net_0[12]\, DRAM_DQ_OE(11) => 
        \DRAM_DQ_OE_net_0[11]\, DRAM_DQ_OE(10) => 
        \DRAM_DQ_OE_net_0[10]\, DRAM_DQ_OE(9) => 
        \DRAM_DQ_OE_net_0[9]\, DRAM_DQ_OE(8) => 
        \DRAM_DQ_OE_net_0[8]\, DRAM_DQ_OE(7) => 
        \DRAM_DQ_OE_net_0[7]\, DRAM_DQ_OE(6) => 
        \DRAM_DQ_OE_net_0[6]\, DRAM_DQ_OE(5) => 
        \DRAM_DQ_OE_net_0[5]\, DRAM_DQ_OE(4) => 
        \DRAM_DQ_OE_net_0[4]\, DRAM_DQ_OE(3) => 
        \DRAM_DQ_OE_net_0[3]\, DRAM_DQ_OE(2) => 
        \DRAM_DQ_OE_net_0[2]\, DRAM_DQ_OE(1) => 
        \DRAM_DQ_OE_net_0[1]\, DRAM_DQ_OE(0) => 
        \DRAM_DQ_OE_net_0[0]\, DRAM_DQS_OE(2) => nc123, 
        DRAM_DQS_OE(1) => \DRAM_DQS_OE_net_0[1]\, DRAM_DQS_OE(0)
         => \DRAM_DQS_OE_net_0[0]\, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, SPI1_SCK_OE => 
        OPEN, SPI1_SDI_MGPIO11A_OE => OPEN, SPI1_SDO_MGPIO12A_OE
         => OPEN, SPI1_SS0_MGPIO13A_OE => OPEN, 
        SPI1_SS1_MGPIO14A_OE => OPEN, SPI1_SS2_MGPIO15A_OE => 
        OPEN, SPI1_SS3_MGPIO16A_OE => OPEN, SPI1_SS4_MGPIO17A_OE
         => OPEN, SPI1_SS5_MGPIO18A_OE => OPEN, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN);
    
    MDDR_RAS_N_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_RASN, PAD => MDDR_RAS_N);
    
    MSS_ADLIB_INST_RNIHJLG_15 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[16]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(16));
    
    MDDR_DQ_4_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(4), D => \DRAM_DQ_OUT_net_0[4]\, E
         => \DRAM_DQ_OE_net_0[4]\, Y => MDDR_DQ_4_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_6 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[7]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(7));
    
    MSS_ADLIB_INST_RNIHJLG_18 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[19]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(19));
    
    MDDR_ADDR_10_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[10]\, PAD => MDDR_ADDR(10));
    
    MDDR_DQS_TMATCH_0_IN_PAD : INBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQS_TMATCH_0_IN, Y => 
        MDDR_DQS_TMATCH_0_IN_PAD_Y);
    
    MDDR_CS_N_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CSN, PAD => MDDR_CS_N);
    
    MSS_ADLIB_INST_RNIHJLG_25 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[26]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(26));
    
    MDDR_ADDR_4_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[4]\, PAD => MDDR_ADDR(4));
    
    MSS_ADLIB_INST_RNIHJLG_28 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[29]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(29));
    
    MDDR_DQ_7_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(7), D => \DRAM_DQ_OUT_net_0[7]\, E
         => \DRAM_DQ_OE_net_0[7]\, Y => MDDR_DQ_7_PAD_Y);
    
    MDDR_WE_N_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_WEN, PAD => MDDR_WE_N);
    
    MSS_ADLIB_INST_RNIHJLG_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[1]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(1));
    
    MSS_ADLIB_INST_RNIHJLG_4 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[5]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(5));
    
    MDDR_ADDR_8_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[8]\, PAD => MDDR_ADDR(8));
    
    MDDR_ADDR_15_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[15]\, PAD => MDDR_ADDR(15));
    
    MDDR_ADDR_0_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[0]\, PAD => MDDR_ADDR(0));
    
    MDDR_ADDR_1_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[1]\, PAD => MDDR_ADDR(1));
    
    MSS_ADLIB_INST_RNIHJLG_10 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[11]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(11));
    
    MSS_ADLIB_INST_RNIHJLG_30 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[31]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(31));
    
    MSS_ADLIB_INST_RNIHJLG_12 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[13]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(13));
    
    MDDR_DQ_13_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(13), D => \DRAM_DQ_OUT_net_0[13]\, 
        E => \DRAM_DQ_OE_net_0[13]\, Y => MDDR_DQ_13_PAD_Y);
    
    MDDR_ADDR_3_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_ADDR_net_0[3]\, PAD => MDDR_ADDR(3));
    
    MSS_ADLIB_INST_RNI67N2 : CLKINT
      port map(A => CONFIG_PRESET_N, Y => 
        \CORECONFIGP_0_APB_S_PRESET_N\);
    
    MDDR_BA_0_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_BA_net_0[0]\, PAD => MDDR_BA(0));
    
    MDDR_DQ_6_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(6), D => \DRAM_DQ_OUT_net_0[6]\, E
         => \DRAM_DQ_OE_net_0[6]\, Y => MDDR_DQ_6_PAD_Y);
    
    MDDR_CLK_PAD : OUTBUF_DIFF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CLK, PADP => MDDR_CLK, 
        PADN => MDDR_CLK_N);
    
    MDDR_DQ_14_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(14), D => \DRAM_DQ_OUT_net_0[14]\, 
        E => \DRAM_DQ_OE_net_0[14]\, Y => MDDR_DQ_14_PAD_Y);
    
    MSS_ADLIB_INST_RNIHJLG_20 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[21]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(21));
    
    MSS_ADLIB_INST_RNIHJLG_22 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[23]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(23));
    
    MSS_ADLIB_INST_RNIHJLG_1 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[2]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(2));
    
    MDDR_DQS_TMATCH_0_OUT_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_FIFO_WE_OUT_net_0[0]\, PAD => 
        MDDR_DQS_TMATCH_0_OUT);
    
    MSS_ADLIB_INST_RNIHJLG_3 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[4]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(4));
    
    MDDR_BA_1_PAD : OUTBUF
      generic map(IOSTD => "LPDDRI")

      port map(D => \DRAM_BA_net_0[1]\, PAD => MDDR_BA(1));
    
    MSS_ADLIB_INST_RNIHJLG_19 : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[20]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(20));
    
    MSS_ADLIB_INST_RNIHJLG : CFG2
      generic map(INIT => x"8")

      port map(A => \CoreAHBLite_1_AHBmslave16_HRDATA[0]\, B => 
        xhdl1328_i_m_0_1(0), Y => ConfigMaster_0_M_HRDATA(0));
    
    MDDR_DQ_5_PAD : BIBUF
      generic map(IOSTD => "LPDDRI")

      port map(PAD => MDDR_DQ(5), D => \DRAM_DQ_OUT_net_0[5]\, E
         => \DRAM_DQ_OE_net_0[5]\, Y => MDDR_DQ_5_PAD_Y);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIU0V1 : CLKINT
      port map(A => FIC_2_APB_M_PCLK, Y => 
        \CORECONFIGP_0_APB_S_PCLK\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Igloo2_TFT_Video_Out_Test_CCC_0_FCCC is

    port( Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0            : out   std_logic;
          HPMS_DDR_FIC_SUBSYSTEM_LOCK                        : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic
        );

end Igloo2_TFT_Video_Out_Test_CCC_0_FCCC;

architecture DEF_ARCH of Igloo2_TFT_Video_Out_Test_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044D64000F18C2718C231839DEC0404041000301",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK, BUSY => OPEN, CLK0 => 
        VCC_net_1, CLK1 => VCC_net_1, CLK2 => VCC_net_1, CLK3 => 
        VCC_net_1, NGMUX0_SEL => GND_net_1, NGMUX1_SEL => 
        GND_net_1, NGMUX2_SEL => GND_net_1, NGMUX3_SEL => 
        GND_net_1, NGMUX0_HOLD_N => VCC_net_1, NGMUX1_HOLD_N => 
        VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, NGMUX3_HOLD_N => 
        VCC_net_1, NGMUX0_ARST_N => VCC_net_1, NGMUX1_ARST_N => 
        VCC_net_1, NGMUX2_ARST_N => VCC_net_1, NGMUX3_ARST_N => 
        VCC_net_1, PLL_BYPASS_N => VCC_net_1, PLL_ARST_N => 
        VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, GPD0_ARST_N => 
        VCC_net_1, GPD1_ARST_N => VCC_net_1, GPD2_ARST_N => 
        VCC_net_1, GPD3_ARST_N => VCC_net_1, PRESET_N => 
        GND_net_1, PCLK => VCC_net_1, PSEL => VCC_net_1, PENABLE
         => VCC_net_1, PWRITE => VCC_net_1, PADDR(7) => VCC_net_1, 
        PADDR(6) => VCC_net_1, PADDR(5) => VCC_net_1, PADDR(4)
         => VCC_net_1, PADDR(3) => VCC_net_1, PADDR(2) => 
        VCC_net_1, PWDATA(7) => VCC_net_1, PWDATA(6) => VCC_net_1, 
        PWDATA(5) => VCC_net_1, PWDATA(4) => VCC_net_1, PWDATA(3)
         => VCC_net_1, PWDATA(2) => VCC_net_1, PWDATA(1) => 
        VCC_net_1, PWDATA(0) => VCC_net_1, CLK0_PAD => GND_net_1, 
        CLK1_PAD => GND_net_1, CLK2_PAD => GND_net_1, CLK3_PAD
         => GND_net_1, GL0 => GL0_net, GL1 => OPEN, GL2 => OPEN, 
        GL3 => OPEN, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreConfigP is

    port( Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA    : in    std_logic_vector(16 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA                         : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR                          : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA                         : in    std_logic_vector(15 downto 0);
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11  : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13  : in    std_logic;
          CORECONFIGP_0_SOFT_RESET_F2M_i_0                            : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY    : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                                : in    std_logic;
          CORECONFIGP_0_APB_S_PCLK                                    : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR   : out   std_logic;
          CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET                : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                                  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                                  : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE                         : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE    : in    std_logic;
          CORECONFIGP_0_APB_S_PCLK_i_0                                : in    std_logic;
          INIT_DONE                                                   : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE                        : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE   : in    std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx     : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx                          : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR                        : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY                         : in    std_logic
        );

end CoreConfigP;

architecture DEF_ARCH of CoreConfigP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal CORECONFIGP_0_SOFT_RESET_F2M, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY\, 
        GND_net_1, \FIC_2_APB_M_PREADY_0_ldmx\, N_52_i_0, 
        VCC_net_1, \prdata[0]\, \state[1]_net_1\, \prdata[1]\, 
        \prdata[2]\, \prdata[3]\, \prdata[4]\, \prdata[5]\, 
        \prdata[6]\, \prdata[7]\, \prdata[8]\, \prdata[9]\, 
        \prdata[10]\, \prdata[11]\, \prdata[12]\, \prdata[13]\, 
        \prdata[14]\, \prdata[15]\, N_27_i_0, N_29_i_0, pslverr, 
        \soft_reset_reg[0]_net_1\, \un17_int_psel_0_a4\, 
        \soft_reset_reg[2]_net_1\, 
        \CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET\, 
        \soft_reset_reg[4]_net_1\, \soft_reset_reg[5]_net_1\, 
        \soft_reset_reg[6]_net_1\, \soft_reset_reg[7]_net_1\, 
        \soft_reset_reg[8]_net_1\, \soft_reset_reg[9]_net_1\, 
        \soft_reset_reg[10]_net_1\, \soft_reset_reg[11]_net_1\, 
        \soft_reset_reg[12]_net_1\, \soft_reset_reg[13]_net_1\, 
        \soft_reset_reg[14]_net_1\, \soft_reset_reg[15]_net_1\, 
        \soft_reset_reg[16]_net_1\, \CORECONFIGP_0_CONFIG1_DONE\, 
        \control_reg_1_ldmx[0]_net_1\, \psel\, 
        \CORECONFIGP_0_CONFIG2_DONE\, 
        \control_reg_1_ldmx[1]_net_1\, \state_d[2]\, 
        \paddr[12]_net_1\, \paddr[13]_net_1\, \paddr[15]_net_1\, 
        \state[0]_net_1\, \state_ns[0]\, \state_ns[1]\, 
        \state_d_i_0[2]\, \INIT_DONE_q1\, \INIT_DONE_q2\, 
        MDDR_PENABLE_0_1, \prdata_0_iv_0_a4_0[12]\, 
        \prdata_0_iv_0_a4_0[9]\, \prdata_0_iv_0_a4_0[10]\, 
        \prdata_0_iv_0_a4_0[15]\, \prdata_0_iv_0_a4_0[7]\, 
        \prdata_0_iv_0_a4_0[8]\, \prdata_0_iv_0_a4_0[2]\, 
        \prdata_0_iv_0_a4_0[4]\, \prdata_0_iv_0_a4_0[11]\, 
        \prdata_0_iv_0_a4_0[14]\, \prdata_0_iv_0_a4_0[13]\, 
        \prdata_0_iv_0_a4_0[3]\, \prdata_0_iv_0_a4_0[6]\, N_92, 
        N_91, N_80, N_43, \control_reg_1_en_2[0]_net_1\, N_44, 
        N_99, \prdata_0_iv_0_a4_1[0]\, \un17_int_psel_0_a4_2\, 
        \un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_a4_0_1\, 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, 
        \control_reg_1_en_4[0]_net_1\, 
        \prdata_0_iv_0_0_a1[5]_net_1\, 
        \prdata_0_iv_0_0_a0[0]_net_1\, 
        \prdata_0_iv_0_0_a0[1]_net_1\ : std_logic;

begin 

    Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY <= 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY\;
    CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET <= 
        \CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET\;
    CORECONFIGP_0_CONFIG1_DONE <= \CORECONFIGP_0_CONFIG1_DONE\;
    CORECONFIGP_0_CONFIG2_DONE <= \CORECONFIGP_0_CONFIG2_DONE\;
    CORECONFIGP_0_MDDR_APBmslave_PSELx <= 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\;

    \soft_reset_reg[13]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(13), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[13]_net_1\);
    
    \pwdata[15]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(15), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15));
    
    \prdata_0_iv_0[1]\ : CFG4
      generic map(INIT => x"F111")

      port map(A => N_99, B => \prdata_0_iv_0_0_a0[1]_net_1\, C
         => CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[1]\);
    
    \pwdata[8]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(8), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8));
    
    \prdata_0_iv_i_a4[16]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \soft_reset_reg[16]_net_1\, B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        Y => N_80);
    
    \pwdata[3]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(3), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3));
    
    \prdata_0_iv_0[15]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), C => 
        \prdata_0_iv_0_a4_0[15]\, D => N_99, Y => \prdata[15]\);
    
    \soft_reset_reg[10]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(10), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[10]_net_1\);
    
    \paddr[8]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8));
    
    \soft_reset_reg[2]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(2), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[2]_net_1\);
    
    \pwdata[5]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(5), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5));
    
    \state_ns_0_0[1]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \state[0]_net_1\, B => 
        \un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_a4_0_1\, C => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, Y => \state_ns[1]\);
    
    \prdata_0_iv_0_a4_0_0[15]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[15]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[15]\);
    
    \paddr[5]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5));
    
    \prdata_0_iv_0_a4_0_0[12]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[12]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[12]\);
    
    INIT_DONE_q1 : SLE
      port map(D => INIT_DONE, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \INIT_DONE_q1\);
    
    \FIC_2_APB_M_PRDATA_0[7]\ : SLE
      port map(D => \prdata[7]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7);
    
    \paddr[3]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3));
    
    \control_reg_1_en_4[0]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        C => \paddr[13]_net_1\, D => 
        \control_reg_1_en_2[0]_net_1\, Y => 
        \control_reg_1_en_4[0]_net_1\);
    
    \pwdata[9]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(9), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9));
    
    \control_reg_1[0]\ : SLE
      port map(D => \control_reg_1_ldmx[0]_net_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \psel\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG1_DONE\);
    
    \pwdata[7]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(7), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7));
    
    FIC_2_APB_M_PREADY_0 : SLE
      port map(D => \FIC_2_APB_M_PREADY_0_ldmx\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => N_52_i_0, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY\);
    
    \soft_reset_reg[9]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(9), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[9]_net_1\);
    
    \control_reg_1_ldmx[1]\ : CFG4
      generic map(INIT => x"E2F0")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(1), 
        B => \paddr[15]_net_1\, C => \CORECONFIGP_0_CONFIG2_DONE\, 
        D => \control_reg_1_en_4[0]_net_1\, Y => 
        \control_reg_1_ldmx[1]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \pwdata[1]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(1), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1));
    
    \pwdata[13]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(13), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13));
    
    \FIC_2_APB_M_PRDATA_0_RNO[16]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        C => N_99, D => N_80, Y => N_27_i_0);
    
    psel : SLE
      port map(D => \state_d_i_0[2]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i_0, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => \psel\);
    
    \FIC_2_APB_M_PRDATA_0[17]\ : SLE
      port map(D => N_29_i_0, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state[1]_net_1\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18);
    
    \FIC_2_APB_M_PRDATA_0[14]\ : SLE
      port map(D => \prdata[14]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14);
    
    pwrite : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE);
    
    \pwdata[6]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(6), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6));
    
    \prdata_0_iv_0_a4_1_0[0]\ : CFG3
      generic map(INIT => x"04")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => N_43, C => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_1[0]\);
    
    \paddr[12]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \paddr[12]_net_1\);
    
    MDDR_PENABLE_0_1_0_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => \paddr[15]_net_1\, B => \paddr[12]_net_1\, Y
         => N_91);
    
    \control_reg_1_en_2[0]\ : CFG3
      generic map(INIT => x"02")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        C => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        Y => \control_reg_1_en_2[0]_net_1\);
    
    \prdata_0_iv_0_a4_0_0[2]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[2]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[2]\);
    
    \paddr[13]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \paddr[13]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[1]\ : SLE
      port map(D => \prdata[1]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1);
    
    un8_int_psel_0_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        Y => N_92);
    
    \soft_reset_reg[0]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(0), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[0]_net_1\);
    
    \pwdata[2]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(2), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2));
    
    \soft_reset_reg_RNIIT9F[1]\ : CFG1
      generic map(INIT => "01")

      port map(A => CORECONFIGP_0_SOFT_RESET_F2M, Y => 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0);
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_o3 : CFG3
      generic map(INIT => x"FD")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        C => \state[0]_net_1\, Y => N_44);
    
    \prdata_0_iv_0_a4_0_0[10]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[10]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[10]\);
    
    \FIC_2_APB_M_PRDATA_0[9]\ : SLE
      port map(D => \prdata[9]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9);
    
    \prdata_0_iv_0_0_a0[5]\ : CFG3
      generic map(INIT => x"C4")

      port map(A => \paddr[13]_net_1\, B => \psel\, C => 
        \paddr[15]_net_1\, Y => N_99);
    
    \FIC_2_APB_M_PRDATA_0[13]\ : SLE
      port map(D => \prdata[13]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13);
    
    \soft_reset_reg[15]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(15), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[15]_net_1\);
    
    \paddr[7]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7));
    
    \FIC_2_APB_M_PRDATA_0[11]\ : SLE
      port map(D => \prdata[11]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11);
    
    \prdata_0_iv_0[9]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), C => 
        \prdata_0_iv_0_a4_0[9]\, D => N_99, Y => \prdata[9]\);
    
    \prdata_0_iv_0_a4_0_0[8]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[8]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[8]\);
    
    \prdata_0_iv_0[7]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), C => 
        \prdata_0_iv_0_a4_0[7]\, D => N_99, Y => \prdata[7]\);
    
    \prdata_0_iv_0_a4_0_0[11]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[11]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[11]\);
    
    \prdata_0_iv_0[0]\ : CFG4
      generic map(INIT => x"F111")

      port map(A => N_99, B => \prdata_0_iv_0_0_a0[0]_net_1\, C
         => CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[0]\);
    
    \paddr[6]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6));
    
    \control_reg_1[1]\ : SLE
      port map(D => \control_reg_1_ldmx[1]_net_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \psel\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG2_DONE\);
    
    \pwdata[11]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(11), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11));
    
    \prdata_0_iv_0[13]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), C => 
        \prdata_0_iv_0_a4_0[13]\, D => N_99, Y => \prdata[13]\);
    
    \FIC_2_APB_M_PRDATA_0[2]\ : SLE
      port map(D => \prdata[2]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \prdata_0_iv_0[14]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), C => 
        \prdata_0_iv_0_a4_0[14]\, D => N_99, Y => \prdata[14]\);
    
    \soft_reset_reg[3]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(3), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        \CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET\);
    
    \soft_reset_reg[12]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(12), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[12]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[8]\ : SLE
      port map(D => \prdata[8]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8);
    
    \state[0]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[0]_net_1\);
    
    \prdata_0_iv_0_0_a0[1]\ : CFG4
      generic map(INIT => x"5D7F")

      port map(A => N_92, B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        C => CORECONFIGP_0_SOFT_RESET_F2M, D => 
        \CORECONFIGP_0_CONFIG2_DONE\, Y => 
        \prdata_0_iv_0_0_a0[1]_net_1\);
    
    state_s0_0_a2_0_a4 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d[2]\);
    
    \prdata_0_iv_0_a4_0_0[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[4]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[4]\);
    
    \prdata_0_iv_0[8]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), C => 
        \prdata_0_iv_0_a4_0[8]\, D => N_99, Y => \prdata[8]\);
    
    \prdata_0_iv_0[10]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), C => 
        \prdata_0_iv_0_a4_0[10]\, D => N_99, Y => \prdata[10]\);
    
    \prdata_0_iv_0_a4_0_0[14]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[14]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[14]\);
    
    \prdata_0_iv_0[6]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), C => 
        \prdata_0_iv_0_a4_0[6]\, D => N_99, Y => \prdata[6]\);
    
    \FIC_2_APB_M_PRDATA_0[10]\ : SLE
      port map(D => \prdata[10]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10);
    
    \pwdata[14]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(14), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14));
    
    \FIC_2_APB_M_PRDATA_0[16]\ : SLE
      port map(D => N_27_i_0, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state[1]_net_1\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16);
    
    \prdata_0_iv_0_m3[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \CORECONFIGP_0_CONFIG1_DONE\, B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \INIT_DONE_q2\, Y => N_43);
    
    FIC_2_APB_M_PREADY_0_ldmx : CFG3
      generic map(INIT => x"EA")

      port map(A => \state[1]_net_1\, B => N_44, C => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY\, 
        Y => \FIC_2_APB_M_PREADY_0_ldmx\);
    
    \soft_reset_reg[4]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(4), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[4]_net_1\);
    
    FIC_2_APB_M_PSLVERR_0 : SLE
      port map(D => pslverr, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state[1]_net_1\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR);
    
    \soft_reset_reg[8]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(8), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[8]_net_1\);
    
    FIC_2_APB_M_PREADY_0_RNO : CFG2
      generic map(INIT => x"B")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PREADY, B => 
        \un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_a4_0_1\, Y => 
        N_52_i_0);
    
    \FIC_2_APB_M_PRDATA_0[3]\ : SLE
      port map(D => \prdata[3]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3);
    
    \prdata_0_iv_0_a4_0_0[6]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[6]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[6]\);
    
    MDDR_PSEL_0_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => \psel\, B => \paddr[13]_net_1\, C => N_91, Y
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\);
    
    un17_int_psel_0_a4 : CFG4
      generic map(INIT => x"4000")

      port map(A => \paddr[15]_net_1\, B => 
        \un17_int_psel_0_a4_2\, C => \psel\, D => 
        \paddr[13]_net_1\, Y => \un17_int_psel_0_a4\);
    
    \pwdata[10]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(10), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10));
    
    INIT_DONE_q2 : SLE
      port map(D => \INIT_DONE_q1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INIT_DONE_q2\);
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_a4_0_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => \state[1]_net_1\, B => \paddr[13]_net_1\, C
         => \psel\, D => N_91, Y => 
        \un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_i_a4_0_1\);
    
    \prdata_0_iv_0[11]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), C => 
        \prdata_0_iv_0_a4_0[11]\, D => N_99, Y => \prdata[11]\);
    
    \FIC_2_APB_M_PRDATA_0[0]\ : SLE
      port map(D => \prdata[0]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0);
    
    \state[1]\ : SLE
      port map(D => \state_ns[1]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[1]_net_1\);
    
    \soft_reset_reg[6]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(6), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[6]_net_1\);
    
    \prdata_0_iv_0[3]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), C => 
        \prdata_0_iv_0_a4_0[3]\, D => N_99, Y => \prdata[3]\);
    
    \prdata_0_iv_0_a4_0_0[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET\, D
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[3]\);
    
    FIC_2_APB_M_PSLVERR_0_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PSLVERR, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => pslverr);
    
    un17_int_psel_0_a4_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_92, B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        C => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \un17_int_psel_0_a4_2\);
    
    \soft_reset_reg[7]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(7), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[7]_net_1\);
    
    \soft_reset_reg[11]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(11), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[11]_net_1\);
    
    \paddr[4]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4));
    
    MDDR_PENABLE_0_1_0_a4 : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[15]_net_1\, C
         => \paddr[13]_net_1\, D => \state[1]_net_1\, Y => 
        MDDR_PENABLE_0_1);
    
    \pwdata[12]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(12), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12));
    
    \paddr[9]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9));
    
    \FIC_2_APB_M_PRDATA_0[15]\ : SLE
      port map(D => \prdata[15]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15);
    
    \soft_reset_reg[1]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(1), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => CORECONFIGP_0_SOFT_RESET_F2M);
    
    \prdata_0_iv_0_a4_0_0[13]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[13]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[13]\);
    
    \soft_reset_reg[16]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(16), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[16]_net_1\);
    
    \pwdata[0]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(0), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0));
    
    \FIC_2_APB_M_PRDATA_0[4]\ : SLE
      port map(D => \prdata[4]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4);
    
    \pwdata[4]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(4), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4));
    
    MDDR_PENABLE_0 : SLE
      port map(D => MDDR_PENABLE_0_1, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i_0, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE);
    
    \prdata_0_iv_0[2]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), C => 
        \prdata_0_iv_0_a4_0[2]\, D => N_99, Y => \prdata[2]\);
    
    \FIC_2_APB_M_PRDATA_0[12]\ : SLE
      port map(D => \prdata[12]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12);
    
    \prdata_0_iv_0_a4_0_0[9]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[9]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[9]\);
    
    \prdata_0_iv_0_0_a1[5]\ : CFG4
      generic map(INIT => x"BDBF")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        C => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        D => \soft_reset_reg[5]_net_1\, Y => 
        \prdata_0_iv_0_0_a1[5]_net_1\);
    
    \prdata_0_iv_0[12]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), C => 
        \prdata_0_iv_0_a4_0[12]\, D => N_99, Y => \prdata[12]\);
    
    \paddr[2]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2));
    
    \prdata_0_iv_0_a4_0_0[7]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        C => \soft_reset_reg[7]_net_1\, D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        Y => \prdata_0_iv_0_a4_0[7]\);
    
    \paddr[10]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10));
    
    psel_RNO : CFG2
      generic map(INIT => x"E")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d_i_0[2]\);
    
    \control_reg_1_ldmx[0]\ : CFG4
      generic map(INIT => x"E2F0")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(0), 
        B => \paddr[15]_net_1\, C => \CORECONFIGP_0_CONFIG1_DONE\, 
        D => \control_reg_1_en_4[0]_net_1\, Y => 
        \control_reg_1_ldmx[0]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[6]\ : SLE
      port map(D => \prdata[6]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6);
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_a3_0_a4 : CFG2
      generic map(INIT => x"1")

      port map(A => N_44, B => \state[1]_net_1\, Y => 
        \state_ns[0]\);
    
    \prdata_0_iv_0[5]\ : CFG4
      generic map(INIT => x"F111")

      port map(A => N_99, B => \prdata_0_iv_0_0_a1[5]_net_1\, C
         => CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[5]\);
    
    \prdata_0_iv_0[4]\ : CFG4
      generic map(INIT => x"88F8")

      port map(A => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), C => 
        \prdata_0_iv_0_a4_0[4]\, D => N_99, Y => \prdata[4]\);
    
    \FIC_2_APB_M_PRDATA_0_RNO[17]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0, 
        B => N_99, C => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1, 
        Y => N_29_i_0);
    
    \soft_reset_reg[14]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(14), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[14]_net_1\);
    
    \prdata_0_iv_0_0_a0[0]\ : CFG4
      generic map(INIT => x"007F")

      port map(A => N_92, B => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2, 
        C => \soft_reset_reg[0]_net_1\, D => 
        \prdata_0_iv_0_a4_1[0]\, Y => 
        \prdata_0_iv_0_0_a0[0]_net_1\);
    
    \paddr[15]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13, 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \paddr[15]_net_1\);
    
    \soft_reset_reg[5]\ : SLE
      port map(D => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(5), 
        CLK => CORECONFIGP_0_APB_S_PCLK, EN => 
        \un17_int_psel_0_a4\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \soft_reset_reg[5]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[5]\ : SLE
      port map(D => \prdata[5]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1 is

    port( xhdl1222                                : in    std_logic_vector(16 to 16);
          SDATASELInt_fast_14                     : in    std_logic;
          SDATASELInt_fast_4                      : in    std_logic;
          SDATASELInt_fast_2                      : in    std_logic;
          SDATASELInt_fast_0                      : in    std_logic;
          SDATASELInt_fast_13                     : in    std_logic;
          SDATASELInt_fast_12                     : in    std_logic;
          SDATASELInt_fast_11                     : in    std_logic;
          SDATASELInt_fast_10                     : in    std_logic;
          SDATASELInt_10                          : in    std_logic;
          SDATASELInt_14                          : in    std_logic;
          SDATASELInt_4                           : in    std_logic;
          SDATASELInt_2                           : in    std_logic;
          SDATASELInt_0                           : in    std_logic;
          SDATASELInt_9                           : in    std_logic;
          SDATASELInt_8                           : in    std_logic;
          SDATASELInt_7                           : in    std_logic;
          SDATASELInt_6                           : in    std_logic;
          SDATASELInt_13                          : in    std_logic;
          SDATASELInt_12                          : in    std_logic;
          SDATASELInt_11                          : in    std_logic;
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          N_107                                   : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          N_106                                   : out   std_logic;
          N_108                                   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic;
          PREVDATASLAVEREADY_iv_i_0               : out   std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1;

architecture DEF_ARCH of 
        COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \defSlaveSMCurrentState\, VCC_net_1, N_4_i_0, 
        GND_net_1, \defSlaveSMNextState_m_0_2_a1_x_sx\, 
        \defSlaveSMNextState_m_0_2_a1_0\, 
        \defSlaveSMNextState_i_a2_0_x\, 
        defSlaveSMNextState_m_0_4_1, 
        \defSlaveSMNextState_m_0_2_a0_x_sx_0\, 
        \defSlaveSMNextState_m_0_2_a0_x_sx\, 
        \defSlaveSMCurrentState_RNISA5T3\, N_112, \N_107\, 
        \defSlaveSMNextState_m_0_2\, 
        \defSlaveSMNextState_m_0_a7_0_0\, 
        \defSlaveSMNextState_m_0_2_a0_0\, 
        \defSlaveSMNextState_m_0_a7_3_0\, \N_106\, \N_108\, 
        \defSlaveSMNextState_m_0_3_1_tz_tz\, \N_98\, \N_25\, 
        \defSlaveSMNextState_m_0_3_1\, 
        \defSlaveSMNextState_m_0_3\ : std_logic;

begin 

    N_107 <= \N_107\;
    defSlaveSMNextState_m_0_2 <= \defSlaveSMNextState_m_0_2\;
    N_106 <= \N_106\;
    N_108 <= \N_108\;
    N_98 <= \N_98\;
    N_25 <= \N_25\;
    defSlaveSMNextState_m_0_3_1 <= \defSlaveSMNextState_m_0_3_1\;
    defSlaveSMNextState_m_0_3 <= \defSlaveSMNextState_m_0_3\;

    defSlaveSMCurrentState : SLE
      port map(D => N_4_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \defSlaveSMCurrentState\);
    
    defSlaveSMNextState_i_a2_0_RNI7CIMC : CFG3
      generic map(INIT => x"FE")

      port map(A => \N_98\, B => \N_25\, C => 
        \defSlaveSMNextState_m_0_3_1\, Y => 
        \defSlaveSMNextState_m_0_3\);
    
    defSlaveSMNextState_m_0_2_a1_0 : CFG4
      generic map(INIT => x"0110")

      port map(A => SDATASELInt_9, B => SDATASELInt_8, C => 
        SDATASELInt_7, D => SDATASELInt_6, Y => 
        \defSlaveSMNextState_m_0_2_a1_0\);
    
    defSlaveSMCurrentState_RNO : CFG4
      generic map(INIT => x"1333")

      port map(A => \N_106\, B => \defSlaveSMCurrentState\, C => 
        \N_107\, D => \N_108\, Y => N_4_i_0);
    
    defSlaveSMCurrentState_RNISA5T3 : CFG4
      generic map(INIT => x"0001")

      port map(A => \defSlaveSMNextState_m_0_2_a0_x_sx_0\, B => 
        \defSlaveSMNextState_m_0_2_a0_x_sx\, C => 
        \defSlaveSMCurrentState\, D => xhdl1222(16), Y => 
        \defSlaveSMCurrentState_RNISA5T3\);
    
    defSlaveSMCurrentState_RNII1HGN : CFG3
      generic map(INIT => x"01")

      port map(A => \defSlaveSMNextState_m_0_3\, B => 
        un1_state_31_i_i_a2_0_d_1_0_1, C => 
        \defSlaveSMNextState_m_0_2\, Y => HREADY_i_3_i_0);
    
    defSlaveSMNextState_m_0_3_1_tz_tz : CFG4
      generic map(INIT => x"0116")

      port map(A => SDATASELInt_13, B => SDATASELInt_12, C => 
        SDATASELInt_11, D => SDATASELInt_10, Y => 
        \defSlaveSMNextState_m_0_3_1_tz_tz\);
    
    defSlaveSMNextState_i_a2_0_x : CFG3
      generic map(INIT => x"01")

      port map(A => SDATASELInt_fast_13, B => SDATASELInt_fast_12, 
        C => SDATASELInt_fast_11, Y => 
        \defSlaveSMNextState_i_a2_0_x\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    defSlaveSMNextState_m_0_2_a0_x_sx_0 : CFG4
      generic map(INIT => x"FFEB")

      port map(A => SDATASELInt_fast_14, B => SDATASELInt_fast_4, 
        C => SDATASELInt_fast_2, D => SDATASELInt_fast_0, Y => 
        \defSlaveSMNextState_m_0_2_a0_x_sx_0\);
    
    defSlaveSMNextState_i_a2_0_RNI9U9KM : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \N_98\, B => \N_25\, C => 
        \defSlaveSMNextState_m_0_3_1\, D => 
        \defSlaveSMNextState_m_0_2\, Y => defSlaveSMNextState_m);
    
    \defSlaveSMNextState_i_a2_0_RNI3J724_1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_106\, B => \N_108\, C => N_112, D => 
        \defSlaveSMNextState_m_0_2_a1_0\, Y => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1);
    
    defSlaveSMNextState_m_0_a2_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_9, B => SDATASELInt_8, C => 
        SDATASELInt_7, D => SDATASELInt_6, Y => \N_107\);
    
    \defSlaveSMNextState_i_a2_0_RNI3J724_2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_108\, B => \N_107\, C => N_112, D => 
        \defSlaveSMNextState_m_0_2_a0_0\, Y => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2);
    
    defSlaveSMCurrentState_RNIQHV4N : CFG3
      generic map(INIT => x"01")

      port map(A => \defSlaveSMNextState_m_0_2\, B => 
        \defSlaveSMNextState_m_0_3\, C => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, Y => 
        PREVDATASLAVEREADY_iv_i_0);
    
    defSlaveSMNextState_m_0_a7_3_0 : CFG4
      generic map(INIT => x"0006")

      port map(A => SDATASELInt_9, B => SDATASELInt_8, C => 
        SDATASELInt_7, D => SDATASELInt_6, Y => 
        \defSlaveSMNextState_m_0_a7_3_0\);
    
    defSlaveSMNextState_m_0_2_a0_0 : CFG4
      generic map(INIT => x"0014")

      port map(A => SDATASELInt_14, B => SDATASELInt_4, C => 
        SDATASELInt_2, D => SDATASELInt_0, Y => 
        \defSlaveSMNextState_m_0_2_a0_0\);
    
    defSlaveSMNextState_i_a2_0_RNI3J724_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_106\, B => \N_108\, C => N_112, D => 
        \defSlaveSMNextState_m_0_a7_3_0\, Y => \N_98\);
    
    defSlaveSMNextState_i_a2_0_RNI3J724 : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_108\, B => \N_107\, C => N_112, D => 
        \defSlaveSMNextState_m_0_a7_0_0\, Y => \N_25\);
    
    defSlaveSMNextState_i_a2_0 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_13, B => SDATASELInt_12, C => 
        SDATASELInt_11, D => SDATASELInt_10, Y => \N_108\);
    
    defSlaveSMNextState_m_0_a7_0_0 : CFG4
      generic map(INIT => x"0102")

      port map(A => SDATASELInt_14, B => SDATASELInt_4, C => 
        SDATASELInt_2, D => SDATASELInt_0, Y => 
        \defSlaveSMNextState_m_0_a7_0_0\);
    
    defSlaveSMNextState_m_0_a2_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => SDATASELInt_14, B => SDATASELInt_4, C => 
        SDATASELInt_2, D => SDATASELInt_0, Y => \N_106\);
    
    defSlaveSMCurrentState_RNI2INT9 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \defSlaveSMCurrentState_RNISA5T3\, B => 
        defSlaveSMNextState_m_0_4_1, C => N_112, D => \N_107\, Y
         => \defSlaveSMNextState_m_0_2\);
    
    defSlaveSMNextState_m_0_2_a0_x_sx : CFG4
      generic map(INIT => x"FFFE")

      port map(A => SDATASELInt_fast_12, B => SDATASELInt_fast_11, 
        C => SDATASELInt_fast_10, D => SDATASELInt_fast_13, Y => 
        \defSlaveSMNextState_m_0_2_a0_x_sx\);
    
    defSlaveSMCurrentState_RNI163I4 : CFG4
      generic map(INIT => x"8000")

      port map(A => \N_106\, B => \N_107\, C => N_112, D => 
        \defSlaveSMNextState_m_0_3_1_tz_tz\, Y => 
        \defSlaveSMNextState_m_0_3_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    defSlaveSMNextState_i_a2_0_x_RNIQ56T3 : CFG4
      generic map(INIT => x"0400")

      port map(A => \defSlaveSMNextState_m_0_2_a1_x_sx\, B => 
        \defSlaveSMNextState_m_0_2_a1_0\, C => SDATASELInt_10, D
         => \defSlaveSMNextState_i_a2_0_x\, Y => 
        defSlaveSMNextState_m_0_4_1);
    
    defSlaveSMNextState_m_0_2_a1_x_sx : CFG4
      generic map(INIT => x"FFFE")

      port map(A => SDATASELInt_fast_14, B => SDATASELInt_fast_4, 
        C => SDATASELInt_fast_2, D => SDATASELInt_fast_0, Y => 
        \defSlaveSMNextState_m_0_2_a1_x_sx\);
    
    defSlaveSMCurrentState_RNIV9TD : CFG2
      generic map(INIT => x"1")

      port map(A => xhdl1222(16), B => \defSlaveSMCurrentState\, 
        Y => N_112);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_1_1_85_65536 is

    port( regHSIZE                                : out   std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0);
          xhdl1222                                : out   std_logic_vector(16 to 16);
          xhdl1221                                : out   std_logic_vector(16 to 16);
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0);
          M0GATEDHADDR                            : out   std_logic_vector(31 downto 29);
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1);
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          regHADDR_0                              : out   std_logic;
          regHADDR_1                              : out   std_logic;
          regHADDR_2                              : out   std_logic;
          regHADDR_3                              : out   std_logic;
          regHADDR_4                              : out   std_logic;
          regHADDR_5                              : out   std_logic;
          regHADDR_6                              : out   std_logic;
          regHADDR_7                              : out   std_logic;
          regHADDR_8                              : out   std_logic;
          regHADDR_9                              : out   std_logic;
          regHADDR_10                             : out   std_logic;
          regHADDR_11                             : out   std_logic;
          regHADDR_12                             : out   std_logic;
          regHADDR_13                             : out   std_logic;
          regHADDR_14                             : out   std_logic;
          regHADDR_15                             : out   std_logic;
          regHADDR_16                             : out   std_logic;
          regHADDR_17                             : out   std_logic;
          regHADDR_18                             : out   std_logic;
          regHADDR_19                             : out   std_logic;
          regHADDR_20                             : out   std_logic;
          regHADDR_21                             : out   std_logic;
          regHADDR_22                             : out   std_logic;
          regHADDR_23                             : out   std_logic;
          regHADDR_24                             : out   std_logic;
          regHADDR_25                             : out   std_logic;
          regHADDR_26                             : out   std_logic;
          regHADDR_27                             : out   std_logic;
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          regHWRITE                               : out   std_logic;
          ConfigMaster_0_M_HWRITE                 : in    std_logic;
          masterRegAddrSel                        : out   std_logic;
          M0GATEDHTRANS                           : out   std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_m      : in    std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic
        );

end COREAHBLITE_MASTERSTAGE_1_1_85_65536;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_1_1_85_65536 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1
    port( xhdl1222                                : in    std_logic_vector(16 to 16) := (others => 'U');
          SDATASELInt_fast_14                     : in    std_logic := 'U';
          SDATASELInt_fast_4                      : in    std_logic := 'U';
          SDATASELInt_fast_2                      : in    std_logic := 'U';
          SDATASELInt_fast_0                      : in    std_logic := 'U';
          SDATASELInt_fast_13                     : in    std_logic := 'U';
          SDATASELInt_fast_12                     : in    std_logic := 'U';
          SDATASELInt_fast_11                     : in    std_logic := 'U';
          SDATASELInt_fast_10                     : in    std_logic := 'U';
          SDATASELInt_10                          : in    std_logic := 'U';
          SDATASELInt_14                          : in    std_logic := 'U';
          SDATASELInt_4                           : in    std_logic := 'U';
          SDATASELInt_2                           : in    std_logic := 'U';
          SDATASELInt_0                           : in    std_logic := 'U';
          SDATASELInt_9                           : in    std_logic := 'U';
          SDATASELInt_8                           : in    std_logic := 'U';
          SDATASELInt_7                           : in    std_logic := 'U';
          SDATASELInt_6                           : in    std_logic := 'U';
          SDATASELInt_13                          : in    std_logic := 'U';
          SDATASELInt_12                          : in    std_logic := 'U';
          SDATASELInt_11                          : in    std_logic := 'U';
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          N_107                                   : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          N_106                                   : out   std_logic;
          N_108                                   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic := 'U';
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic := 'U';
          PREVDATASLAVEREADY_iv_i_0               : out   std_logic
        );
  end component;

    signal VCC_net_1, \masterAddrClockEnable\, GND_net_1, 
        \regHADDR[29]_net_1\, \regHADDR[30]_net_1\, \regHTRANS\, 
        \SDATASELInt[1]_net_1\, \SADDRSEL[1]_net_1\, 
        PREVDATASLAVEREADY_iv_i_0, \SDATASELInt[3]_net_1\, 
        \SADDRSEL[3]_net_1\, \SDATASELInt[5]_net_1\, 
        \SADDRSEL[5]_net_1\, \SDATASELInt[7]_net_1\, 
        \SADDRSEL[7]_net_1\, \SDATASELInt[8]_net_1\, 
        \SADDRSEL[8]_net_1\, \SDATASELInt[9]_net_1\, 
        \SADDRSEL[9]_net_1\, \SDATASELInt[10]_net_1\, 
        \SADDRSEL[10]_net_1\, \SDATASELInt[11]_net_1\, 
        \SADDRSEL[11]_net_1\, \SDATASELInt[12]_net_1\, 
        \SADDRSEL[12]_net_1\, \SDATASELInt[13]_net_1\, 
        \SADDRSEL[13]_net_1\, \SDATASELInt[14]_net_1\, 
        \SADDRSEL[14]_net_1\, \SDATASELInt[15]_net_1\, 
        \SADDRSEL[15]_net_1\, \xhdl1222[16]\, \xhdl1221[16]\, 
        masterRegAddrSel_net_1, \d_masterRegAddrSel\, 
        \SDATASELInt_fast[15]_net_1\, \SADDRSEL_fast[15]_net_1\, 
        \SDATASELInt_fast[1]_net_1\, \SADDRSEL_fast[1]_net_1\, 
        \SDATASELInt_fast[3]_net_1\, \SADDRSEL_fast[3]_net_1\, 
        \SDATASELInt_fast[5]_net_1\, \SADDRSEL_fast[5]_net_1\, 
        \SDATASELInt_fast[12]_net_1\, \SADDRSEL_fast[12]_net_1\, 
        \SDATASELInt_fast[14]_net_1\, \SADDRSEL_fast[14]_net_1\, 
        \SDATASELInt_fast[13]_net_1\, \SADDRSEL_fast[13]_net_1\, 
        \SDATASELInt_fast[11]_net_1\, \SADDRSEL_fast[11]_net_1\, 
        \M0GATEDHTRANS\, \M0GATEDHADDR[31]\, \M0GATEDHADDR[30]\, 
        \SADDRSEL_1[7]\, \M0GATEDHADDR[29]\, 
        \SADDRSEL_0[14]_net_1\, \SADDRSEL_2[12]\, 
        \SADDRSEL_0[8]_net_1\, N_106, N_107, N_108, 
        \defSlaveSMNextState_m_0_3\, \defSlaveSMNextState_m_0_2\, 
        \HREADY_i_3\ : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1
	Use entity work.
        COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1(DEF_ARCH);
begin 

    xhdl1222(16) <= \xhdl1222[16]\;
    xhdl1221(16) <= \xhdl1221[16]\;
    M0GATEDHADDR(31) <= \M0GATEDHADDR[31]\;
    M0GATEDHADDR(30) <= \M0GATEDHADDR[30]\;
    M0GATEDHADDR(29) <= \M0GATEDHADDR[29]\;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    M0GATEDHTRANS <= \M0GATEDHTRANS\;
    defSlaveSMNextState_m_0_3 <= \defSlaveSMNextState_m_0_3\;
    defSlaveSMNextState_m_0_2 <= \defSlaveSMNextState_m_0_2\;
    HREADY_i_3 <= \HREADY_i_3\;

    \SADDRSEL[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => ConfigMaster_0_M_HADDR(30), B => 
        \M0GATEDHTRANS\, C => \M0GATEDHADDR[29]\, D => 
        \SADDRSEL_2[12]\, Y => \SADDRSEL[12]_net_1\);
    
    \regHADDR[21]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(21), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_21);
    
    \PREGATEDHADDR[31]\ : CFG2
      generic map(INIT => x"4")

      port map(A => masterRegAddrSel_net_1, B => 
        ConfigMaster_0_M_HADDR(31), Y => \M0GATEDHADDR[31]\);
    
    \regHADDR[15]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(15), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_15);
    
    \SADDRSEL[13]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[13]_net_1\);
    
    \regHADDR[30]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(30), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \regHADDR[30]_net_1\);
    
    \regHADDR[7]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(7), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_7);
    
    \SADDRSEL_fast[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[3]_net_1\);
    
    \SADDRSEL[1]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => ConfigMaster_0_M_HADDR(29), B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[31]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[1]_net_1\);
    
    \SADDRSEL[9]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => ConfigMaster_0_M_HADDR(31), B => 
        ConfigMaster_0_M_HADDR(29), C => \SADDRSEL_1[7]\, D => 
        \M0GATEDHADDR[30]\, Y => \SADDRSEL[9]_net_1\);
    
    \SADDRSEL[16]\ : CFG4
      generic map(INIT => x"F010")

      port map(A => ConfigMaster_0_M_HADDR(28), B => 
        ConfigMaster_0_M_HADDR(31), C => \M0GATEDHTRANS\, D => 
        masterRegAddrSel_net_1, Y => \xhdl1221[16]\);
    
    \PREGATEDHADDR[30]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[30]_net_1\, B => 
        masterRegAddrSel_net_1, C => ConfigMaster_0_M_HADDR(30), 
        Y => \M0GATEDHADDR[30]\);
    
    \regHADDR[9]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(9), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_9);
    
    \SADDRSEL[11]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(29), C => \M0GATEDHADDR[30]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[11]_net_1\);
    
    \masterRegAddrSel\ : SLE
      port map(D => \d_masterRegAddrSel\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        masterRegAddrSel_net_1);
    
    regHTRANS : SLE
      port map(D => VCC_net_1, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \regHTRANS\);
    
    \SDATASELInt_fast[14]\ : SLE
      port map(D => \SADDRSEL_fast[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[14]_net_1\);
    
    GATEDHTRANS : CFG3
      generic map(INIT => x"D8")

      port map(A => masterRegAddrSel_net_1, B => \regHTRANS\, C
         => ConfigMaster_0_M_HTRANS(1), Y => \M0GATEDHTRANS\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \SADDRSEL_fast[13]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[13]_net_1\);
    
    \SADDRSEL_fast[5]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[5]_net_1\);
    
    \regHADDR[29]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(29), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \regHADDR[29]_net_1\);
    
    \SADDRSEL_fast[15]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => ConfigMaster_0_M_HADDR(29), B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[31]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[15]_net_1\);
    
    \SADDRSEL_fast[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \M0GATEDHADDR[29]\, B => 
        \SADDRSEL_0[14]_net_1\, C => \M0GATEDHTRANS\, Y => 
        \SADDRSEL_fast[14]_net_1\);
    
    \SADDRSEL_1[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ConfigMaster_0_M_HADDR(28), B => 
        masterRegAddrSel_net_1, C => ConfigMaster_0_M_HTRANS(1), 
        Y => \SADDRSEL_1[7]\);
    
    \SADDRSEL[15]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => ConfigMaster_0_M_HADDR(29), B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[31]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[15]_net_1\);
    
    \regHADDR[24]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(24), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_24);
    
    \SDATASELInt_fast[11]\ : SLE
      port map(D => \SADDRSEL_fast[11]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[11]_net_1\);
    
    \regHADDR[10]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(10), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_10);
    
    \regHADDR[13]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(13), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_13);
    
    \regHADDR[12]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(12), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_12);
    
    \regHADDR[5]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(5), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_5);
    
    \SADDRSEL[8]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \SADDRSEL_0[8]_net_1\, B => 
        \M0GATEDHADDR[31]\, C => \M0GATEDHADDR[30]\, D => 
        \M0GATEDHADDR[29]\, Y => \SADDRSEL[8]_net_1\);
    
    \regHADDR[2]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(2), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_2);
    
    \SDATASELInt[15]\ : SLE
      port map(D => \SADDRSEL[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[15]_net_1\);
    
    \SADDRSEL[10]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \M0GATEDHADDR[29]\, B => \SADDRSEL_2[12]\, C
         => \M0GATEDHTRANS\, D => \M0GATEDHADDR[30]\, Y => 
        \SADDRSEL[10]_net_1\);
    
    \SDATASELInt[14]\ : SLE
      port map(D => \SADDRSEL[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[14]_net_1\);
    
    \regHADDR[8]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(8), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_8);
    
    \regHADDR[25]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(25), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_25);
    
    \SDATASELInt_fast[3]\ : SLE
      port map(D => \SADDRSEL_fast[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[3]_net_1\);
    
    \SDATASELInt_fast[13]\ : SLE
      port map(D => \SADDRSEL_fast[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[13]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SADDRSEL_fast[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => ConfigMaster_0_M_HADDR(30), B => 
        \M0GATEDHTRANS\, C => \M0GATEDHADDR[29]\, D => 
        \SADDRSEL_2[12]\, Y => \SADDRSEL_fast[12]_net_1\);
    
    \SADDRSEL_0[8]\ : CFG3
      generic map(INIT => x"D0")

      port map(A => ConfigMaster_0_M_HADDR(28), B => 
        masterRegAddrSel_net_1, C => ConfigMaster_0_M_HTRANS(1), 
        Y => \SADDRSEL_0[8]_net_1\);
    
    \regHADDR[17]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(17), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_17);
    
    \SDATASELInt_fast[12]\ : SLE
      port map(D => \SADDRSEL_fast[12]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[12]_net_1\);
    
    \SADDRSEL[7]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => ConfigMaster_0_M_HADDR(29), B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[31]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[7]_net_1\);
    
    masterAddrClockEnable : CFG4
      generic map(INIT => x"0100")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY_m, B => 
        \HREADY_i_3\, C => masterRegAddrSel_net_1, D => 
        \xhdl1221[16]\, Y => \masterAddrClockEnable\);
    
    \SDATASELInt_fast[15]\ : SLE
      port map(D => \SADDRSEL_fast[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[15]_net_1\);
    
    \regHADDR[6]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(6), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_6);
    
    \regHADDR[16]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(16), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_16);
    
    \SDATASELInt[13]\ : SLE
      port map(D => \SADDRSEL[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[13]_net_1\);
    
    \regHWRITE\ : SLE
      port map(D => ConfigMaster_0_M_HWRITE, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHWRITE);
    
    \regHSIZE[1]\ : SLE
      port map(D => ConfigMaster_0_M_HSIZE(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHSIZE(1));
    
    d_masterRegAddrSel : CFG4
      generic map(INIT => x"5100")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY_m, B => 
        \HREADY_i_3\, C => masterRegAddrSel_net_1, D => 
        \xhdl1221[16]\, Y => \d_masterRegAddrSel\);
    
    \SDATASELInt[9]\ : SLE
      port map(D => \SADDRSEL[9]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[9]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => \SADDRSEL[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[1]_net_1\);
    
    \SDATASELInt[12]\ : SLE
      port map(D => \SADDRSEL[12]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[12]_net_1\);
    
    \SADDRSEL_fast[1]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => ConfigMaster_0_M_HADDR(29), B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[31]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[1]_net_1\);
    
    \regHADDR[11]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(11), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_11);
    
    \regHADDR[0]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_0);
    
    HREADY_M_iv : CFG3
      generic map(INIT => x"FE")

      port map(A => \defSlaveSMNextState_m_0_3\, B => 
        un1_state_31_i_i_a2_0_d_1_0_1, C => 
        \defSlaveSMNextState_m_0_2\, Y => \HREADY_i_3\);
    
    \SADDRSEL[5]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[5]_net_1\);
    
    \SDATASELInt[5]\ : SLE
      port map(D => \SADDRSEL[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[5]_net_1\);
    
    \regHADDR[3]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(3), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_3);
    
    \SADDRSEL[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \M0GATEDHADDR[29]\, B => 
        \SADDRSEL_0[14]_net_1\, C => \M0GATEDHTRANS\, Y => 
        \SADDRSEL[14]_net_1\);
    
    \SDATASELInt[3]\ : SLE
      port map(D => \SADDRSEL[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[3]_net_1\);
    
    \SADDRSEL_fast[11]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(29), C => \M0GATEDHADDR[30]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL_fast[11]_net_1\);
    
    \regHADDR[20]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(20), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_20);
    
    \regHADDR[23]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(23), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_23);
    
    \regHADDR[1]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_1);
    
    \regHADDR[22]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(22), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_22);
    
    \SDATASELInt[7]\ : SLE
      port map(D => \SADDRSEL[7]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[7]_net_1\);
    
    \regHSIZE[0]\ : SLE
      port map(D => ConfigMaster_0_M_HSIZE(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHSIZE(0));
    
    hready_m_xhdl355_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_106, B => \xhdl1222[16]\, C => N_107, D => 
        N_108, Y => xhdl1328_i_m_0_1(0));
    
    \SADDRSEL_2[10]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(28), Y => \SADDRSEL_2[12]\);
    
    \PREGATEDHADDR[29]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \regHADDR[29]_net_1\, B => 
        masterRegAddrSel_net_1, C => ConfigMaster_0_M_HADDR(29), 
        Y => \M0GATEDHADDR[29]\);
    
    \regHADDR[19]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(19), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_19);
    
    \regHADDR[14]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(14), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_14);
    
    \regHADDR[27]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(27), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_27);
    
    \SDATASELInt[16]\ : SLE
      port map(D => \xhdl1221[16]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \xhdl1222[16]\);
    
    \SADDRSEL[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \M0GATEDHADDR[31]\, B => 
        ConfigMaster_0_M_HADDR(30), C => \M0GATEDHADDR[29]\, D
         => \SADDRSEL_1[7]\, Y => \SADDRSEL[3]_net_1\);
    
    \regHADDR[18]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(18), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_18);
    
    \SDATASELInt[11]\ : SLE
      port map(D => \SADDRSEL[11]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[11]_net_1\);
    
    \SDATASELInt_fast[1]\ : SLE
      port map(D => \SADDRSEL_fast[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[1]_net_1\);
    
    \SDATASELInt[8]\ : SLE
      port map(D => \SADDRSEL[8]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[8]_net_1\);
    
    \SADDRSEL_0[14]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => ConfigMaster_0_M_HADDR(31), B => 
        ConfigMaster_0_M_HADDR(28), C => masterRegAddrSel_net_1, 
        D => ConfigMaster_0_M_HADDR(30), Y => 
        \SADDRSEL_0[14]_net_1\);
    
    \regHADDR[4]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(4), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_4);
    
    \regHADDR[26]\ : SLE
      port map(D => ConfigMaster_0_M_HADDR(26), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \masterAddrClockEnable\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => regHADDR_26);
    
    \SDATASELInt[10]\ : SLE
      port map(D => \SADDRSEL[10]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[10]_net_1\);
    
    \SDATASELInt_fast[5]\ : SLE
      port map(D => \SADDRSEL_fast[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        PREVDATASLAVEREADY_iv_i_0, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt_fast[5]_net_1\);
    
    default_slave_sm : 
        COREAHBLITE_DEFAULTSLAVESM_default_slave_sm_1
      port map(xhdl1222(16) => \xhdl1222[16]\, 
        SDATASELInt_fast_14 => \SDATASELInt_fast[15]_net_1\, 
        SDATASELInt_fast_4 => \SDATASELInt_fast[5]_net_1\, 
        SDATASELInt_fast_2 => \SDATASELInt_fast[3]_net_1\, 
        SDATASELInt_fast_0 => \SDATASELInt_fast[1]_net_1\, 
        SDATASELInt_fast_13 => \SDATASELInt_fast[14]_net_1\, 
        SDATASELInt_fast_12 => \SDATASELInt_fast[13]_net_1\, 
        SDATASELInt_fast_11 => \SDATASELInt_fast[12]_net_1\, 
        SDATASELInt_fast_10 => \SDATASELInt_fast[11]_net_1\, 
        SDATASELInt_10 => \SDATASELInt[11]_net_1\, SDATASELInt_14
         => \SDATASELInt[15]_net_1\, SDATASELInt_4 => 
        \SDATASELInt[5]_net_1\, SDATASELInt_2 => 
        \SDATASELInt[3]_net_1\, SDATASELInt_0 => 
        \SDATASELInt[1]_net_1\, SDATASELInt_9 => 
        \SDATASELInt[10]_net_1\, SDATASELInt_8 => 
        \SDATASELInt[9]_net_1\, SDATASELInt_7 => 
        \SDATASELInt[8]_net_1\, SDATASELInt_6 => 
        \SDATASELInt[7]_net_1\, SDATASELInt_13 => 
        \SDATASELInt[14]_net_1\, SDATASELInt_12 => 
        \SDATASELInt[13]_net_1\, SDATASELInt_11 => 
        \SDATASELInt[12]_net_1\, HPMS_READY => HPMS_READY, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, N_107 => N_107, 
        defSlaveSMNextState_m_0_2 => \defSlaveSMNextState_m_0_2\, 
        N_106 => N_106, N_108 => N_108, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, N_98 => N_98, N_25
         => N_25, defSlaveSMNextState_m_0_3_1 => 
        defSlaveSMNextState_m_0_3_1, defSlaveSMNextState_m_0_3
         => \defSlaveSMNextState_m_0_3\, defSlaveSMNextState_m
         => defSlaveSMNextState_m, un1_state_31_i_i_a2_0_d_1_0_1
         => un1_state_31_i_i_a2_0_d_1_0_1, HREADY_i_3_i_0 => 
        HREADY_i_3_i_0, CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, 
        PREVDATASLAVEREADY_iv_i_0 => PREVDATASLAVEREADY_iv_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_slave_arbiter_2 is

    port( masterAddrInProg                        : out   std_logic_vector(3 downto 1);
          xhdl1221                                : in    std_logic_vector(16 to 16);
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic;
          N_152                                   : out   std_logic;
          N_152_i_0                               : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_m      : out   std_logic
        );

end COREAHBLITE_SLAVEARBITER_slave_arbiter_2;

architecture DEF_ARCH of 
        COREAHBLITE_SLAVEARBITER_slave_arbiter_2 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[1]_net_1\, VCC_net_1, N_126_i_0, 
        GND_net_1, \masterAddrInProg[3]\, N_128_i_0, 
        \arbRegSMCurrentState[15]_net_1\, N_104_i_0, 
        \arbRegSMCurrentState[14]_net_1\, N_106_i_0, 
        \arbRegSMCurrentState[13]_net_1\, N_108_i_0, 
        \arbRegSMCurrentState[12]_net_1\, N_110_i_0, 
        \arbRegSMCurrentState[10]_net_1\, 
        \arbRegSMCurrentState_ns[5]_net_1\, 
        \arbRegSMCurrentState[9]_net_1\, N_114_i_0, 
        \masterAddrInProg[1]\, N_116_i_0, 
        \arbRegSMCurrentState[6]_net_1\, 
        \arbRegSMCurrentState_ns[9]_net_1\, 
        \arbRegSMCurrentState[5]_net_1\, N_120_i_0, 
        \masterAddrInProg[2]\, N_122_i_0, 
        \arbRegSMCurrentState[2]_net_1\, 
        \arbRegSMCurrentState_ns[13]_net_1\, N_106_i_1, N_139, 
        N_156, \N_152\ : std_logic;

begin 

    masterAddrInProg(3) <= \masterAddrInProg[3]\;
    masterAddrInProg(2) <= \masterAddrInProg[2]\;
    masterAddrInProg(1) <= \masterAddrInProg[1]\;
    N_152 <= \N_152\;

    \arbRegSMCurrentState_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[3]\, Y => N_126_i_0);
    
    \arbRegSMCurrentState_ns_i_a2_0_RNIPATV[0]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => N_156, B => xhdl1221(16), C => 
        \arbRegSMCurrentState[15]_net_1\, D => 
        \arbRegSMCurrentState[12]_net_1\, Y => N_152_i_0);
    
    \arbRegSMCurrentState_ns[13]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[1]_net_1\, B => 
        \arbRegSMCurrentState[2]_net_1\, C => xhdl1221(16), Y => 
        \arbRegSMCurrentState_ns[13]_net_1\);
    
    \arbRegSMCurrentState[12]\ : SLE
      port map(D => N_110_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[12]_net_1\);
    
    \arbRegSMCurrentState_ns[9]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[5]_net_1\, B => 
        \arbRegSMCurrentState[6]_net_1\, C => xhdl1221(16), Y => 
        \arbRegSMCurrentState_ns[9]_net_1\);
    
    \arbRegSMCurrentState[8]\ : SLE
      port map(D => N_116_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[1]\);
    
    \arbRegSMCurrentState[10]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[10]_net_1\);
    
    \arbRegSMCurrentState_RNO_0[14]\ : CFG4
      generic map(INIT => x"1151")

      port map(A => \arbRegSMCurrentState[13]_net_1\, B => 
        \arbRegSMCurrentState[14]_net_1\, C => xhdl1221(16), D
         => CoreAHBLite_1_AHBmslave16_HREADY, Y => N_106_i_1);
    
    \MASTERADDRINPROG_i_a2[0]\ : CFG4
      generic map(INIT => x"000B")

      port map(A => N_156, B => xhdl1221(16), C => 
        \arbRegSMCurrentState[15]_net_1\, D => 
        \arbRegSMCurrentState[12]_net_1\, Y => \N_152\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[3]\, Y => N_128_i_0);
    
    \arbRegSMCurrentState[0]\ : SLE
      port map(D => N_128_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[3]\);
    
    \arbRegSMCurrentState_RNO[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \arbRegSMCurrentState[12]_net_1\, Y => N_110_i_0);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG4
      generic map(INIT => x"0D0C")

      port map(A => N_156, B => \arbRegSMCurrentState[15]_net_1\, 
        C => CoreAHBLite_1_AHBmslave16_HREADY, D => xhdl1221(16), 
        Y => N_104_i_0);
    
    \arbRegSMCurrentState_RNO[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[1]\, Y => N_116_i_0);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_106_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[14]_net_1\);
    
    \arbRegSMCurrentState_ns_i_o2_0[1]\ : CFG4
      generic map(INIT => x"3337")

      port map(A => \arbRegSMCurrentState[2]_net_1\, B => 
        xhdl1221(16), C => \arbRegSMCurrentState[10]_net_1\, D
         => \arbRegSMCurrentState[6]_net_1\, Y => N_139);
    
    \arbRegSMCurrentState[6]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[9]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[6]_net_1\);
    
    \arbRegSMCurrentState[1]\ : SLE
      port map(D => N_126_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_RNO[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[2]\, Y => N_122_i_0);
    
    \arbRegSMCurrentState_RNO[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \arbRegSMCurrentState[12]_net_1\, Y => N_108_i_0);
    
    \arbRegSMCurrentState_RNO[14]\ : CFG4
      generic map(INIT => x"B3BB")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        N_106_i_1, C => \arbRegSMCurrentState[15]_net_1\, D => 
        N_139, Y => N_106_i_0);
    
    \arbRegSMCurrentState[9]\ : SLE
      port map(D => N_114_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[9]_net_1\);
    
    \arbRegSMCurrentState[4]\ : SLE
      port map(D => N_122_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[2]\);
    
    \arbRegSMCurrentState_ns_i_a2_0[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \arbRegSMCurrentState[14]_net_1\, B => 
        \arbRegSMCurrentState[10]_net_1\, C => 
        \arbRegSMCurrentState[6]_net_1\, D => 
        \arbRegSMCurrentState[2]_net_1\, Y => N_156);
    
    \arbRegSMCurrentState[13]\ : SLE
      port map(D => N_108_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[13]_net_1\);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[2]_net_1\);
    
    \arbRegSMCurrentState[5]\ : SLE
      port map(D => N_120_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[5]_net_1\);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_104_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[15]_net_1\);
    
    \MASTERADDRINPROG_i_a2_RNIAHI6[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \N_152\, Y => CoreAHBLite_1_AHBmslave16_HREADY_m);
    
    \arbRegSMCurrentState_ns[5]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[9]_net_1\, B => 
        \arbRegSMCurrentState[10]_net_1\, C => xhdl1221(16), Y
         => \arbRegSMCurrentState_ns[5]_net_1\);
    
    \arbRegSMCurrentState_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[2]\, Y => N_120_i_0);
    
    \arbRegSMCurrentState_RNO[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAHBLite_1_AHBmslave16_HREADY, B => 
        \masterAddrInProg[1]\, Y => N_114_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_slavestage_16 is

    port( ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          xhdl1328_i_m_0_1                        : in    std_logic_vector(0 to 0);
          ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0);
          regHSIZE                                : in    std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          regHADDR                                : in    std_logic_vector(27 downto 0);
          M0GATEDHADDR                            : in    std_logic_vector(31 downto 29);
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(28 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          xhdl1222                                : in    std_logic_vector(16 to 16);
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          xhdl1221                                : in    std_logic_vector(16 to 16);
          masterDataInProg_0                      : out   std_logic;
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          masterRegAddrSel                        : in    std_logic;
          ConfigMaster_0_M_HWRITE                 : in    std_logic;
          regHWRITE                               : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic;
          defSlaveSMNextState_m                   : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic;
          M0GATEDHTRANS                           : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_m      : out   std_logic
        );

end COREAHBLITE_SLAVESTAGE_slavestage_16;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_slavestage_16 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_slave_arbiter_2
    port( masterAddrInProg                        : out   std_logic_vector(3 downto 1);
          xhdl1221                                : in    std_logic_vector(16 to 16) := (others => 'U');
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic := 'U';
          N_152                                   : out   std_logic;
          N_152_i_0                               : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_m      : out   std_logic
        );
  end component;

    signal \masterDataInProg_0\, VCC_net_1, N_152_i_0, GND_net_1, 
        \masterDataInProg[1]_net_1\, \masterAddrInProg[1]\, 
        \masterDataInProg[2]_net_1\, \masterAddrInProg[2]\, 
        \masterDataInProg[3]_net_1\, \masterAddrInProg[3]\, 
        \hwdata10\, N_152, \hsel2\, \un1_htrans_1\ : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_slave_arbiter_2
	Use entity work.
        COREAHBLITE_SLAVEARBITER_slave_arbiter_2(DEF_ARCH);
begin 

    masterDataInProg_0 <= \masterDataInProg_0\;

    \masterDataInProg[3]\ : SLE
      port map(D => \masterAddrInProg[3]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        CoreAHBLite_1_AHBmslave16_HREADY, ALn => HPMS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \masterDataInProg[3]_net_1\);
    
    hsel2_RNITPSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(9), B => regHADDR(9), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(9));
    
    hwdata10_RNIOMRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(16), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(16));
    
    hwdata10_RNI7KCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(6), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(6));
    
    hwdata10_RNILKSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(22), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(22));
    
    hsel2_RNIPLSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(7), B => regHADDR(7), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(7));
    
    hwdata10_RNIANCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(9), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(9));
    
    hwdata10_RNI5ICD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(4), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(4));
    
    hsel2_RNIO3AG : CFG2
      generic map(INIT => x"8")

      port map(A => \hsel2\, B => M0GATEDHADDR(30), Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(30));
    
    hsel2_RNITQGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(27), B => regHADDR(27), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(27));
    
    hwdata10_RNIQORK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(18), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(18));
    
    hsel2_RNIFBSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(2), B => regHADDR(2), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(2));
    
    un1_htrans_1 : CFG4
      generic map(INIT => x"11F1")

      port map(A => defSlaveSMNextState_m, B => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, C => xhdl1222(16), 
        D => N_152, Y => \un1_htrans_1\);
    
    HTRANS : CFG3
      generic map(INIT => x"80")

      port map(A => M0GATEDHTRANS, B => \hsel2\, C => 
        \un1_htrans_1\, Y => CoreAHBLite_1_AHBmslave16_HTRANS(1));
    
    hsel2_RNI0B9G : CFG2
      generic map(INIT => x"8")

      port map(A => \hsel2\, B => M0GATEDHADDR(29), Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(29));
    
    hwdata10_RNI1ECD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(0), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(0));
    
    hsel2_RNIPMGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(25), B => regHADDR(25), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(25));
    
    hsel2_RNINJSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(6), B => regHADDR(6), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(6));
    
    hwdata10_RNIKIRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(12), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(12));
    
    hsel2_RNIROGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(26), B => regHADDR(26), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(26));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    hwdata10_RNIONSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(25), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(25));
    
    hwdata10_RNIJISK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(20), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(20));
    
    HSEL_1 : CFG4
      generic map(INIT => x"0449")

      port map(A => \masterAddrInProg[1]\, B => N_152, C => 
        \masterAddrInProg[3]\, D => \masterAddrInProg[2]\, Y => 
        CoreAHBLite_1_AHBmslave16_HSELx);
    
    hsel2_RNINKGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(24), B => regHADDR(24), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(24));
    
    \masterDataInProg[2]\ : SLE
      port map(D => \masterAddrInProg[2]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        CoreAHBLite_1_AHBmslave16_HREADY, ALn => HPMS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \masterDataInProg[2]_net_1\);
    
    hwdata10_RNINLRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(15), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(15));
    
    hwdata10_RNIJHRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(11), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(11));
    
    hsel2_RNIVQEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(19), B => regHADDR(19), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(19));
    
    hwdata10_RNIIGRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(10), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(10));
    
    hwdata10_RNIRQSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(28), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(28));
    
    hsel2_RNITOEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(18), B => regHADDR(18), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(18));
    
    hsel2_RNIB7SN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(0), B => regHADDR(0), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(0));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \masterDataInProg[1]\ : SLE
      port map(D => \masterAddrInProg[1]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        CoreAHBLite_1_AHBmslave16_HREADY, ALn => HPMS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \masterDataInProg[1]_net_1\);
    
    \masterDataInProg[0]\ : SLE
      port map(D => N_152_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        CoreAHBLite_1_AHBmslave16_HREADY, ALn => HPMS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \masterDataInProg_0\);
    
    hsel2_RNIJFSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(4), B => regHADDR(4), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(4));
    
    hwdata10_RNIMLSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(23), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(23));
    
    hwdata10_RNI9MCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(8), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(8));
    
    hsel2_RNILIGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(23), B => regHADDR(23), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(23));
    
    hwdata10_RNIMKRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(14), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(14));
    
    hwdata10_RNI4HCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(3), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(3));
    
    hsel2_RNIJEEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(13), B => regHADDR(13), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(13));
    
    hsel2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \masterAddrInProg[1]\, B => N_152, C => 
        \masterAddrInProg[3]\, D => \masterAddrInProg[2]\, Y => 
        \hsel2\);
    
    hwdata10_RNIPNRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(17), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(17));
    
    hwdata10_RNIKKTK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(30), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(30));
    
    hsel2_RNIJGGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(22), B => regHADDR(22), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(22));
    
    hsel2_RNINIEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(15), B => regHADDR(15), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(15));
    
    hwdata10_RNILLTK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(31), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(31));
    
    hsel2_RNIP4AG : CFG2
      generic map(INIT => x"8")

      port map(A => \hsel2\, B => M0GATEDHADDR(31), Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(31));
    
    hsel2_RNIHCEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(12), B => regHADDR(12), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(12));
    
    hsel2_RNIFCGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(20), B => regHADDR(20), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(20));
    
    hwdata10_RNINMSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(24), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(24));
    
    hsel2_RNID9SN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(1), B => regHADDR(1), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(1));
    
    hwdata10_RNIRPRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(19), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(19));
    
    hsel2_RNIHDSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(3), B => regHADDR(3), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(3));
    
    hwdata10_RNI3GCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(2), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(2));
    
    hsel2_RNILHSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(5), B => regHADDR(5), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(5));
    
    hsel2_RNIPKEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(16), B => regHADDR(16), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(16));
    
    hwdata10_RNILJRK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(13), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(13));
    
    hsel2_RNIBLT01 : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HSIZE(0), B => regHSIZE(0), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HSIZE(0));
    
    hsel2_RNILGEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(14), B => regHADDR(14), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(14));
    
    hsel2_RNI76FH : CFG3
      generic map(INIT => x"20")

      port map(A => ConfigMaster_0_M_HADDR(28), B => 
        masterRegAddrSel, C => \hsel2\, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(28));
    
    hwdata10_RNI2FCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(1), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(1));
    
    hsel2_RNID8EI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(10), B => regHADDR(10), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(10));
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_slave_arbiter_2
      port map(masterAddrInProg(3) => \masterAddrInProg[3]\, 
        masterAddrInProg(2) => \masterAddrInProg[2]\, 
        masterAddrInProg(1) => \masterAddrInProg[1]\, 
        xhdl1221(16) => xhdl1221(16), HPMS_READY => HPMS_READY, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, N_152 => N_152, 
        N_152_i_0 => N_152_i_0, 
        CoreAHBLite_1_AHBmslave16_HREADY_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_m);
    
    hsel2_RNIRNSN : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(8), B => regHADDR(8), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(8));
    
    hwdata10_RNI8LCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(7), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(7));
    
    hwdata10 : CFG4
      generic map(INIT => x"0100")

      port map(A => \masterDataInProg[3]_net_1\, B => 
        \masterDataInProg[2]_net_1\, C => 
        \masterDataInProg[1]_net_1\, D => \masterDataInProg_0\, Y
         => \hwdata10\);
    
    hsel2_RNIHEGI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(21), B => regHADDR(21), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(21));
    
    hsel2_RNIDNT01 : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HSIZE(1), B => regHSIZE(1), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HSIZE(1));
    
    hsel2_RNIFAEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(11), B => regHADDR(11), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(11));
    
    hwdata10_RNIQPSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(27), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(27));
    
    hwdata10_RNIPOSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(26), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(26));
    
    hsel2_RNIRTT31 : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HWRITE, B => regHWRITE, C
         => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HWRITE);
    
    hwdata10_RNIKJSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(21), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(21));
    
    \masterDataInProg_RNI937S[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \masterDataInProg_0\, B => 
        xhdl1328_i_m_0_1(0), C => 
        CoreAHBLite_1_AHBmslave16_HREADY, Y => 
        un1_state_31_i_i_a2_0_d_1_0_1);
    
    hwdata10_RNISRSK : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(29), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(29));
    
    hwdata10_RNI6JCD : CFG2
      generic map(INIT => x"8")

      port map(A => \hwdata10\, B => ConfigMaster_0_M_HWDATA(5), 
        Y => CoreAHBLite_1_AHBmslave16_HWDATA(5));
    
    hsel2_RNIRMEI : CFG4
      generic map(INIT => x"C0A0")

      port map(A => ConfigMaster_0_M_HADDR(17), B => regHADDR(17), 
        C => \hsel2\, D => masterRegAddrSel, Y => 
        CoreAHBLite_1_AHBmslave16_HADDR(17));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0 is

    port( ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0);
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1);
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          masterDataInProg                        : out   std_logic_vector(0 to 0);
          ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          ConfigMaster_0_M_HWRITE                 : in    std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic
        );

end COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0;

architecture DEF_ARCH of 
        COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_1_1_85_65536
    port( regHSIZE                                : out   std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          xhdl1222                                : out   std_logic_vector(16 to 16);
          xhdl1221                                : out   std_logic_vector(16 to 16);
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          M0GATEDHADDR                            : out   std_logic_vector(31 downto 29);
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1) := (others => 'U');
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          regHADDR_0                              : out   std_logic;
          regHADDR_1                              : out   std_logic;
          regHADDR_2                              : out   std_logic;
          regHADDR_3                              : out   std_logic;
          regHADDR_4                              : out   std_logic;
          regHADDR_5                              : out   std_logic;
          regHADDR_6                              : out   std_logic;
          regHADDR_7                              : out   std_logic;
          regHADDR_8                              : out   std_logic;
          regHADDR_9                              : out   std_logic;
          regHADDR_10                             : out   std_logic;
          regHADDR_11                             : out   std_logic;
          regHADDR_12                             : out   std_logic;
          regHADDR_13                             : out   std_logic;
          regHADDR_14                             : out   std_logic;
          regHADDR_15                             : out   std_logic;
          regHADDR_16                             : out   std_logic;
          regHADDR_17                             : out   std_logic;
          regHADDR_18                             : out   std_logic;
          regHADDR_19                             : out   std_logic;
          regHADDR_20                             : out   std_logic;
          regHADDR_21                             : out   std_logic;
          regHADDR_22                             : out   std_logic;
          regHADDR_23                             : out   std_logic;
          regHADDR_24                             : out   std_logic;
          regHADDR_25                             : out   std_logic;
          regHADDR_26                             : out   std_logic;
          regHADDR_27                             : out   std_logic;
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          regHWRITE                               : out   std_logic;
          ConfigMaster_0_M_HWRITE                 : in    std_logic := 'U';
          masterRegAddrSel                        : out   std_logic;
          M0GATEDHTRANS                           : out   std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic := 'U';
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_m      : in    std_logic := 'U';
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic := 'U'
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_slavestage_16
    port( ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          xhdl1328_i_m_0_1                        : in    std_logic_vector(0 to 0) := (others => 'U');
          ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          regHSIZE                                : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          regHADDR                                : in    std_logic_vector(27 downto 0) := (others => 'U');
          M0GATEDHADDR                            : in    std_logic_vector(31 downto 29) := (others => 'U');
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(28 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          xhdl1222                                : in    std_logic_vector(16 to 16) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          xhdl1221                                : in    std_logic_vector(16 to 16) := (others => 'U');
          masterDataInProg_0                      : out   std_logic;
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic := 'U';
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          masterRegAddrSel                        : in    std_logic := 'U';
          ConfigMaster_0_M_HWRITE                 : in    std_logic := 'U';
          regHWRITE                               : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic;
          defSlaveSMNextState_m                   : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic := 'U';
          M0GATEDHTRANS                           : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY_m      : out   std_logic
        );
  end component;

    signal \regHADDR[0]\, \regHADDR[1]\, \regHADDR[2]\, 
        \regHADDR[3]\, \regHADDR[4]\, \regHADDR[5]\, 
        \regHADDR[6]\, \regHADDR[7]\, \regHADDR[8]\, 
        \regHADDR[9]\, \regHADDR[10]\, \regHADDR[11]\, 
        \regHADDR[12]\, \regHADDR[13]\, \regHADDR[14]\, 
        \regHADDR[15]\, \regHADDR[16]\, \regHADDR[17]\, 
        \regHADDR[18]\, \regHADDR[19]\, \regHADDR[20]\, 
        \regHADDR[21]\, \regHADDR[22]\, \regHADDR[23]\, 
        \regHADDR[24]\, \regHADDR[25]\, \regHADDR[26]\, 
        \regHADDR[27]\, \regHSIZE[0]\, \regHSIZE[1]\, 
        \xhdl1222[16]\, \xhdl1221[16]\, \M0GATEDHADDR[29]\, 
        \M0GATEDHADDR[30]\, \M0GATEDHADDR[31]\, 
        \xhdl1328_i_m_0_1[0]\, regHWRITE, masterRegAddrSel, 
        M0GATEDHTRANS, \un1_state_31_i_i_a2_0_d_1_0_1\, 
        CoreAHBLite_1_AHBmslave16_HREADY_m, 
        \defSlaveSMNextState_m\, GND_net_1, VCC_net_1
         : std_logic;

    for all : COREAHBLITE_MASTERSTAGE_1_1_85_65536
	Use entity work.COREAHBLITE_MASTERSTAGE_1_1_85_65536(DEF_ARCH);
    for all : COREAHBLITE_SLAVESTAGE_slavestage_16
	Use entity work.COREAHBLITE_SLAVESTAGE_slavestage_16(DEF_ARCH);
begin 

    xhdl1328_i_m_0_1(0) <= \xhdl1328_i_m_0_1[0]\;
    un1_state_31_i_i_a2_0_d_1_0_1 <= 
        \un1_state_31_i_i_a2_0_d_1_0_1\;
    defSlaveSMNextState_m <= \defSlaveSMNextState_m\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_1_1_85_65536
      port map(regHSIZE(1) => \regHSIZE[1]\, regHSIZE(0) => 
        \regHSIZE[0]\, ConfigMaster_0_M_HSIZE(1) => 
        ConfigMaster_0_M_HSIZE(1), ConfigMaster_0_M_HSIZE(0) => 
        ConfigMaster_0_M_HSIZE(0), xhdl1222(16) => \xhdl1222[16]\, 
        xhdl1221(16) => \xhdl1221[16]\, 
        ConfigMaster_0_M_HADDR(31) => ConfigMaster_0_M_HADDR(31), 
        ConfigMaster_0_M_HADDR(30) => ConfigMaster_0_M_HADDR(30), 
        ConfigMaster_0_M_HADDR(29) => ConfigMaster_0_M_HADDR(29), 
        ConfigMaster_0_M_HADDR(28) => ConfigMaster_0_M_HADDR(28), 
        ConfigMaster_0_M_HADDR(27) => ConfigMaster_0_M_HADDR(27), 
        ConfigMaster_0_M_HADDR(26) => ConfigMaster_0_M_HADDR(26), 
        ConfigMaster_0_M_HADDR(25) => ConfigMaster_0_M_HADDR(25), 
        ConfigMaster_0_M_HADDR(24) => ConfigMaster_0_M_HADDR(24), 
        ConfigMaster_0_M_HADDR(23) => ConfigMaster_0_M_HADDR(23), 
        ConfigMaster_0_M_HADDR(22) => ConfigMaster_0_M_HADDR(22), 
        ConfigMaster_0_M_HADDR(21) => ConfigMaster_0_M_HADDR(21), 
        ConfigMaster_0_M_HADDR(20) => ConfigMaster_0_M_HADDR(20), 
        ConfigMaster_0_M_HADDR(19) => ConfigMaster_0_M_HADDR(19), 
        ConfigMaster_0_M_HADDR(18) => ConfigMaster_0_M_HADDR(18), 
        ConfigMaster_0_M_HADDR(17) => ConfigMaster_0_M_HADDR(17), 
        ConfigMaster_0_M_HADDR(16) => ConfigMaster_0_M_HADDR(16), 
        ConfigMaster_0_M_HADDR(15) => ConfigMaster_0_M_HADDR(15), 
        ConfigMaster_0_M_HADDR(14) => ConfigMaster_0_M_HADDR(14), 
        ConfigMaster_0_M_HADDR(13) => ConfigMaster_0_M_HADDR(13), 
        ConfigMaster_0_M_HADDR(12) => ConfigMaster_0_M_HADDR(12), 
        ConfigMaster_0_M_HADDR(11) => ConfigMaster_0_M_HADDR(11), 
        ConfigMaster_0_M_HADDR(10) => ConfigMaster_0_M_HADDR(10), 
        ConfigMaster_0_M_HADDR(9) => ConfigMaster_0_M_HADDR(9), 
        ConfigMaster_0_M_HADDR(8) => ConfigMaster_0_M_HADDR(8), 
        ConfigMaster_0_M_HADDR(7) => ConfigMaster_0_M_HADDR(7), 
        ConfigMaster_0_M_HADDR(6) => ConfigMaster_0_M_HADDR(6), 
        ConfigMaster_0_M_HADDR(5) => ConfigMaster_0_M_HADDR(5), 
        ConfigMaster_0_M_HADDR(4) => ConfigMaster_0_M_HADDR(4), 
        ConfigMaster_0_M_HADDR(3) => ConfigMaster_0_M_HADDR(3), 
        ConfigMaster_0_M_HADDR(2) => ConfigMaster_0_M_HADDR(2), 
        ConfigMaster_0_M_HADDR(1) => ConfigMaster_0_M_HADDR(1), 
        ConfigMaster_0_M_HADDR(0) => ConfigMaster_0_M_HADDR(0), 
        M0GATEDHADDR(31) => \M0GATEDHADDR[31]\, M0GATEDHADDR(30)
         => \M0GATEDHADDR[30]\, M0GATEDHADDR(29) => 
        \M0GATEDHADDR[29]\, ConfigMaster_0_M_HTRANS(1) => 
        ConfigMaster_0_M_HTRANS(1), xhdl1328_i_m_0_1(0) => 
        \xhdl1328_i_m_0_1[0]\, regHADDR_0 => \regHADDR[0]\, 
        regHADDR_1 => \regHADDR[1]\, regHADDR_2 => \regHADDR[2]\, 
        regHADDR_3 => \regHADDR[3]\, regHADDR_4 => \regHADDR[4]\, 
        regHADDR_5 => \regHADDR[5]\, regHADDR_6 => \regHADDR[6]\, 
        regHADDR_7 => \regHADDR[7]\, regHADDR_8 => \regHADDR[8]\, 
        regHADDR_9 => \regHADDR[9]\, regHADDR_10 => 
        \regHADDR[10]\, regHADDR_11 => \regHADDR[11]\, 
        regHADDR_12 => \regHADDR[12]\, regHADDR_13 => 
        \regHADDR[13]\, regHADDR_14 => \regHADDR[14]\, 
        regHADDR_15 => \regHADDR[15]\, regHADDR_16 => 
        \regHADDR[16]\, regHADDR_17 => \regHADDR[17]\, 
        regHADDR_18 => \regHADDR[18]\, regHADDR_19 => 
        \regHADDR[19]\, regHADDR_20 => \regHADDR[20]\, 
        regHADDR_21 => \regHADDR[21]\, regHADDR_22 => 
        \regHADDR[22]\, regHADDR_23 => \regHADDR[23]\, 
        regHADDR_24 => \regHADDR[24]\, regHADDR_25 => 
        \regHADDR[25]\, regHADDR_26 => \regHADDR[26]\, 
        regHADDR_27 => \regHADDR[27]\, HPMS_READY => HPMS_READY, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, regHWRITE => 
        regHWRITE, ConfigMaster_0_M_HWRITE => 
        ConfigMaster_0_M_HWRITE, masterRegAddrSel => 
        masterRegAddrSel, M0GATEDHTRANS => M0GATEDHTRANS, 
        defSlaveSMNextState_m_0_3 => defSlaveSMNextState_m_0_3, 
        un1_state_31_i_i_a2_0_d_1_0_1 => 
        \un1_state_31_i_i_a2_0_d_1_0_1\, 
        defSlaveSMNextState_m_0_2 => defSlaveSMNextState_m_0_2, 
        HREADY_i_3 => HREADY_i_3, 
        CoreAHBLite_1_AHBmslave16_HREADY_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_m, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, N_98 => N_98, N_25
         => N_25, defSlaveSMNextState_m_0_3_1 => 
        defSlaveSMNextState_m_0_3_1, defSlaveSMNextState_m => 
        \defSlaveSMNextState_m\, HREADY_i_3_i_0 => HREADY_i_3_i_0, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m);
    
    slavestage_16 : COREAHBLITE_SLAVESTAGE_slavestage_16
      port map(ConfigMaster_0_M_HWDATA(31) => 
        ConfigMaster_0_M_HWDATA(31), ConfigMaster_0_M_HWDATA(30)
         => ConfigMaster_0_M_HWDATA(30), 
        ConfigMaster_0_M_HWDATA(29) => 
        ConfigMaster_0_M_HWDATA(29), ConfigMaster_0_M_HWDATA(28)
         => ConfigMaster_0_M_HWDATA(28), 
        ConfigMaster_0_M_HWDATA(27) => 
        ConfigMaster_0_M_HWDATA(27), ConfigMaster_0_M_HWDATA(26)
         => ConfigMaster_0_M_HWDATA(26), 
        ConfigMaster_0_M_HWDATA(25) => 
        ConfigMaster_0_M_HWDATA(25), ConfigMaster_0_M_HWDATA(24)
         => ConfigMaster_0_M_HWDATA(24), 
        ConfigMaster_0_M_HWDATA(23) => 
        ConfigMaster_0_M_HWDATA(23), ConfigMaster_0_M_HWDATA(22)
         => ConfigMaster_0_M_HWDATA(22), 
        ConfigMaster_0_M_HWDATA(21) => 
        ConfigMaster_0_M_HWDATA(21), ConfigMaster_0_M_HWDATA(20)
         => ConfigMaster_0_M_HWDATA(20), 
        ConfigMaster_0_M_HWDATA(19) => 
        ConfigMaster_0_M_HWDATA(19), ConfigMaster_0_M_HWDATA(18)
         => ConfigMaster_0_M_HWDATA(18), 
        ConfigMaster_0_M_HWDATA(17) => 
        ConfigMaster_0_M_HWDATA(17), ConfigMaster_0_M_HWDATA(16)
         => ConfigMaster_0_M_HWDATA(16), 
        ConfigMaster_0_M_HWDATA(15) => 
        ConfigMaster_0_M_HWDATA(15), ConfigMaster_0_M_HWDATA(14)
         => ConfigMaster_0_M_HWDATA(14), 
        ConfigMaster_0_M_HWDATA(13) => 
        ConfigMaster_0_M_HWDATA(13), ConfigMaster_0_M_HWDATA(12)
         => ConfigMaster_0_M_HWDATA(12), 
        ConfigMaster_0_M_HWDATA(11) => 
        ConfigMaster_0_M_HWDATA(11), ConfigMaster_0_M_HWDATA(10)
         => ConfigMaster_0_M_HWDATA(10), 
        ConfigMaster_0_M_HWDATA(9) => ConfigMaster_0_M_HWDATA(9), 
        ConfigMaster_0_M_HWDATA(8) => ConfigMaster_0_M_HWDATA(8), 
        ConfigMaster_0_M_HWDATA(7) => ConfigMaster_0_M_HWDATA(7), 
        ConfigMaster_0_M_HWDATA(6) => ConfigMaster_0_M_HWDATA(6), 
        ConfigMaster_0_M_HWDATA(5) => ConfigMaster_0_M_HWDATA(5), 
        ConfigMaster_0_M_HWDATA(4) => ConfigMaster_0_M_HWDATA(4), 
        ConfigMaster_0_M_HWDATA(3) => ConfigMaster_0_M_HWDATA(3), 
        ConfigMaster_0_M_HWDATA(2) => ConfigMaster_0_M_HWDATA(2), 
        ConfigMaster_0_M_HWDATA(1) => ConfigMaster_0_M_HWDATA(1), 
        ConfigMaster_0_M_HWDATA(0) => ConfigMaster_0_M_HWDATA(0), 
        CoreAHBLite_1_AHBmslave16_HWDATA(31) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(31), 
        CoreAHBLite_1_AHBmslave16_HWDATA(30) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(30), 
        CoreAHBLite_1_AHBmslave16_HWDATA(29) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(29), 
        CoreAHBLite_1_AHBmslave16_HWDATA(28) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(28), 
        CoreAHBLite_1_AHBmslave16_HWDATA(27) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(27), 
        CoreAHBLite_1_AHBmslave16_HWDATA(26) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(26), 
        CoreAHBLite_1_AHBmslave16_HWDATA(25) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(25), 
        CoreAHBLite_1_AHBmslave16_HWDATA(24) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(24), 
        CoreAHBLite_1_AHBmslave16_HWDATA(23) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(23), 
        CoreAHBLite_1_AHBmslave16_HWDATA(22) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(22), 
        CoreAHBLite_1_AHBmslave16_HWDATA(21) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(21), 
        CoreAHBLite_1_AHBmslave16_HWDATA(20) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(20), 
        CoreAHBLite_1_AHBmslave16_HWDATA(19) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(19), 
        CoreAHBLite_1_AHBmslave16_HWDATA(18) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(18), 
        CoreAHBLite_1_AHBmslave16_HWDATA(17) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(17), 
        CoreAHBLite_1_AHBmslave16_HWDATA(16) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(16), 
        CoreAHBLite_1_AHBmslave16_HWDATA(15) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(15), 
        CoreAHBLite_1_AHBmslave16_HWDATA(14) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(14), 
        CoreAHBLite_1_AHBmslave16_HWDATA(13) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(13), 
        CoreAHBLite_1_AHBmslave16_HWDATA(12) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(12), 
        CoreAHBLite_1_AHBmslave16_HWDATA(11) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(11), 
        CoreAHBLite_1_AHBmslave16_HWDATA(10) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(10), 
        CoreAHBLite_1_AHBmslave16_HWDATA(9) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(9), 
        CoreAHBLite_1_AHBmslave16_HWDATA(8) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(8), 
        CoreAHBLite_1_AHBmslave16_HWDATA(7) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(7), 
        CoreAHBLite_1_AHBmslave16_HWDATA(6) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(6), 
        CoreAHBLite_1_AHBmslave16_HWDATA(5) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(5), 
        CoreAHBLite_1_AHBmslave16_HWDATA(4) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(4), 
        CoreAHBLite_1_AHBmslave16_HWDATA(3) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(3), 
        CoreAHBLite_1_AHBmslave16_HWDATA(2) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(2), 
        CoreAHBLite_1_AHBmslave16_HWDATA(1) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(1), 
        CoreAHBLite_1_AHBmslave16_HWDATA(0) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(0), xhdl1328_i_m_0_1(0)
         => \xhdl1328_i_m_0_1[0]\, ConfigMaster_0_M_HSIZE(1) => 
        ConfigMaster_0_M_HSIZE(1), ConfigMaster_0_M_HSIZE(0) => 
        ConfigMaster_0_M_HSIZE(0), regHSIZE(1) => \regHSIZE[1]\, 
        regHSIZE(0) => \regHSIZE[0]\, 
        CoreAHBLite_1_AHBmslave16_HSIZE(1) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(1), 
        CoreAHBLite_1_AHBmslave16_HSIZE(0) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(0), regHADDR(27) => 
        \regHADDR[27]\, regHADDR(26) => \regHADDR[26]\, 
        regHADDR(25) => \regHADDR[25]\, regHADDR(24) => 
        \regHADDR[24]\, regHADDR(23) => \regHADDR[23]\, 
        regHADDR(22) => \regHADDR[22]\, regHADDR(21) => 
        \regHADDR[21]\, regHADDR(20) => \regHADDR[20]\, 
        regHADDR(19) => \regHADDR[19]\, regHADDR(18) => 
        \regHADDR[18]\, regHADDR(17) => \regHADDR[17]\, 
        regHADDR(16) => \regHADDR[16]\, regHADDR(15) => 
        \regHADDR[15]\, regHADDR(14) => \regHADDR[14]\, 
        regHADDR(13) => \regHADDR[13]\, regHADDR(12) => 
        \regHADDR[12]\, regHADDR(11) => \regHADDR[11]\, 
        regHADDR(10) => \regHADDR[10]\, regHADDR(9) => 
        \regHADDR[9]\, regHADDR(8) => \regHADDR[8]\, regHADDR(7)
         => \regHADDR[7]\, regHADDR(6) => \regHADDR[6]\, 
        regHADDR(5) => \regHADDR[5]\, regHADDR(4) => 
        \regHADDR[4]\, regHADDR(3) => \regHADDR[3]\, regHADDR(2)
         => \regHADDR[2]\, regHADDR(1) => \regHADDR[1]\, 
        regHADDR(0) => \regHADDR[0]\, M0GATEDHADDR(31) => 
        \M0GATEDHADDR[31]\, M0GATEDHADDR(30) => 
        \M0GATEDHADDR[30]\, M0GATEDHADDR(29) => 
        \M0GATEDHADDR[29]\, ConfigMaster_0_M_HADDR(28) => 
        ConfigMaster_0_M_HADDR(28), ConfigMaster_0_M_HADDR(27)
         => ConfigMaster_0_M_HADDR(27), 
        ConfigMaster_0_M_HADDR(26) => ConfigMaster_0_M_HADDR(26), 
        ConfigMaster_0_M_HADDR(25) => ConfigMaster_0_M_HADDR(25), 
        ConfigMaster_0_M_HADDR(24) => ConfigMaster_0_M_HADDR(24), 
        ConfigMaster_0_M_HADDR(23) => ConfigMaster_0_M_HADDR(23), 
        ConfigMaster_0_M_HADDR(22) => ConfigMaster_0_M_HADDR(22), 
        ConfigMaster_0_M_HADDR(21) => ConfigMaster_0_M_HADDR(21), 
        ConfigMaster_0_M_HADDR(20) => ConfigMaster_0_M_HADDR(20), 
        ConfigMaster_0_M_HADDR(19) => ConfigMaster_0_M_HADDR(19), 
        ConfigMaster_0_M_HADDR(18) => ConfigMaster_0_M_HADDR(18), 
        ConfigMaster_0_M_HADDR(17) => ConfigMaster_0_M_HADDR(17), 
        ConfigMaster_0_M_HADDR(16) => ConfigMaster_0_M_HADDR(16), 
        ConfigMaster_0_M_HADDR(15) => ConfigMaster_0_M_HADDR(15), 
        ConfigMaster_0_M_HADDR(14) => ConfigMaster_0_M_HADDR(14), 
        ConfigMaster_0_M_HADDR(13) => ConfigMaster_0_M_HADDR(13), 
        ConfigMaster_0_M_HADDR(12) => ConfigMaster_0_M_HADDR(12), 
        ConfigMaster_0_M_HADDR(11) => ConfigMaster_0_M_HADDR(11), 
        ConfigMaster_0_M_HADDR(10) => ConfigMaster_0_M_HADDR(10), 
        ConfigMaster_0_M_HADDR(9) => ConfigMaster_0_M_HADDR(9), 
        ConfigMaster_0_M_HADDR(8) => ConfigMaster_0_M_HADDR(8), 
        ConfigMaster_0_M_HADDR(7) => ConfigMaster_0_M_HADDR(7), 
        ConfigMaster_0_M_HADDR(6) => ConfigMaster_0_M_HADDR(6), 
        ConfigMaster_0_M_HADDR(5) => ConfigMaster_0_M_HADDR(5), 
        ConfigMaster_0_M_HADDR(4) => ConfigMaster_0_M_HADDR(4), 
        ConfigMaster_0_M_HADDR(3) => ConfigMaster_0_M_HADDR(3), 
        ConfigMaster_0_M_HADDR(2) => ConfigMaster_0_M_HADDR(2), 
        ConfigMaster_0_M_HADDR(1) => ConfigMaster_0_M_HADDR(1), 
        ConfigMaster_0_M_HADDR(0) => ConfigMaster_0_M_HADDR(0), 
        CoreAHBLite_1_AHBmslave16_HADDR(31) => 
        CoreAHBLite_1_AHBmslave16_HADDR(31), 
        CoreAHBLite_1_AHBmslave16_HADDR(30) => 
        CoreAHBLite_1_AHBmslave16_HADDR(30), 
        CoreAHBLite_1_AHBmslave16_HADDR(29) => 
        CoreAHBLite_1_AHBmslave16_HADDR(29), 
        CoreAHBLite_1_AHBmslave16_HADDR(28) => 
        CoreAHBLite_1_AHBmslave16_HADDR(28), 
        CoreAHBLite_1_AHBmslave16_HADDR(27) => 
        CoreAHBLite_1_AHBmslave16_HADDR(27), 
        CoreAHBLite_1_AHBmslave16_HADDR(26) => 
        CoreAHBLite_1_AHBmslave16_HADDR(26), 
        CoreAHBLite_1_AHBmslave16_HADDR(25) => 
        CoreAHBLite_1_AHBmslave16_HADDR(25), 
        CoreAHBLite_1_AHBmslave16_HADDR(24) => 
        CoreAHBLite_1_AHBmslave16_HADDR(24), 
        CoreAHBLite_1_AHBmslave16_HADDR(23) => 
        CoreAHBLite_1_AHBmslave16_HADDR(23), 
        CoreAHBLite_1_AHBmslave16_HADDR(22) => 
        CoreAHBLite_1_AHBmslave16_HADDR(22), 
        CoreAHBLite_1_AHBmslave16_HADDR(21) => 
        CoreAHBLite_1_AHBmslave16_HADDR(21), 
        CoreAHBLite_1_AHBmslave16_HADDR(20) => 
        CoreAHBLite_1_AHBmslave16_HADDR(20), 
        CoreAHBLite_1_AHBmslave16_HADDR(19) => 
        CoreAHBLite_1_AHBmslave16_HADDR(19), 
        CoreAHBLite_1_AHBmslave16_HADDR(18) => 
        CoreAHBLite_1_AHBmslave16_HADDR(18), 
        CoreAHBLite_1_AHBmslave16_HADDR(17) => 
        CoreAHBLite_1_AHBmslave16_HADDR(17), 
        CoreAHBLite_1_AHBmslave16_HADDR(16) => 
        CoreAHBLite_1_AHBmslave16_HADDR(16), 
        CoreAHBLite_1_AHBmslave16_HADDR(15) => 
        CoreAHBLite_1_AHBmslave16_HADDR(15), 
        CoreAHBLite_1_AHBmslave16_HADDR(14) => 
        CoreAHBLite_1_AHBmslave16_HADDR(14), 
        CoreAHBLite_1_AHBmslave16_HADDR(13) => 
        CoreAHBLite_1_AHBmslave16_HADDR(13), 
        CoreAHBLite_1_AHBmslave16_HADDR(12) => 
        CoreAHBLite_1_AHBmslave16_HADDR(12), 
        CoreAHBLite_1_AHBmslave16_HADDR(11) => 
        CoreAHBLite_1_AHBmslave16_HADDR(11), 
        CoreAHBLite_1_AHBmslave16_HADDR(10) => 
        CoreAHBLite_1_AHBmslave16_HADDR(10), 
        CoreAHBLite_1_AHBmslave16_HADDR(9) => 
        CoreAHBLite_1_AHBmslave16_HADDR(9), 
        CoreAHBLite_1_AHBmslave16_HADDR(8) => 
        CoreAHBLite_1_AHBmslave16_HADDR(8), 
        CoreAHBLite_1_AHBmslave16_HADDR(7) => 
        CoreAHBLite_1_AHBmslave16_HADDR(7), 
        CoreAHBLite_1_AHBmslave16_HADDR(6) => 
        CoreAHBLite_1_AHBmslave16_HADDR(6), 
        CoreAHBLite_1_AHBmslave16_HADDR(5) => 
        CoreAHBLite_1_AHBmslave16_HADDR(5), 
        CoreAHBLite_1_AHBmslave16_HADDR(4) => 
        CoreAHBLite_1_AHBmslave16_HADDR(4), 
        CoreAHBLite_1_AHBmslave16_HADDR(3) => 
        CoreAHBLite_1_AHBmslave16_HADDR(3), 
        CoreAHBLite_1_AHBmslave16_HADDR(2) => 
        CoreAHBLite_1_AHBmslave16_HADDR(2), 
        CoreAHBLite_1_AHBmslave16_HADDR(1) => 
        CoreAHBLite_1_AHBmslave16_HADDR(1), 
        CoreAHBLite_1_AHBmslave16_HADDR(0) => 
        CoreAHBLite_1_AHBmslave16_HADDR(0), xhdl1222(16) => 
        \xhdl1222[16]\, CoreAHBLite_1_AHBmslave16_HTRANS(1) => 
        CoreAHBLite_1_AHBmslave16_HTRANS(1), xhdl1221(16) => 
        \xhdl1221[16]\, masterDataInProg_0 => masterDataInProg(0), 
        HPMS_READY => HPMS_READY, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, 
        un1_state_31_i_i_a2_0_d_1_0_1 => 
        \un1_state_31_i_i_a2_0_d_1_0_1\, 
        CoreAHBLite_1_AHBmslave16_HSELx => 
        CoreAHBLite_1_AHBmslave16_HSELx, masterRegAddrSel => 
        masterRegAddrSel, ConfigMaster_0_M_HWRITE => 
        ConfigMaster_0_M_HWRITE, regHWRITE => regHWRITE, 
        CoreAHBLite_1_AHBmslave16_HWRITE => 
        CoreAHBLite_1_AHBmslave16_HWRITE, defSlaveSMNextState_m
         => \defSlaveSMNextState_m\, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, M0GATEDHTRANS => 
        M0GATEDHTRANS, CoreAHBLite_1_AHBmslave16_HREADY_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_m);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity 
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0 is

    port( ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0);
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1);
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          masterDataInProg                        : out   std_logic_vector(0 to 0);
          ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          ConfigMaster_0_M_HWRITE                 : in    std_logic;
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic
        );

end 
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0;

architecture DEF_ARCH of 
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0
    port( ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1) := (others => 'U');
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          masterDataInProg                        : out   std_logic_vector(0 to 0);
          ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          ConfigMaster_0_M_HWRITE                 : in    std_logic := 'U';
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0
	Use entity work.
        COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0
      port map(ConfigMaster_0_M_HSIZE(1) => 
        ConfigMaster_0_M_HSIZE(1), ConfigMaster_0_M_HSIZE(0) => 
        ConfigMaster_0_M_HSIZE(0), ConfigMaster_0_M_HADDR(31) => 
        ConfigMaster_0_M_HADDR(31), ConfigMaster_0_M_HADDR(30)
         => ConfigMaster_0_M_HADDR(30), 
        ConfigMaster_0_M_HADDR(29) => ConfigMaster_0_M_HADDR(29), 
        ConfigMaster_0_M_HADDR(28) => ConfigMaster_0_M_HADDR(28), 
        ConfigMaster_0_M_HADDR(27) => ConfigMaster_0_M_HADDR(27), 
        ConfigMaster_0_M_HADDR(26) => ConfigMaster_0_M_HADDR(26), 
        ConfigMaster_0_M_HADDR(25) => ConfigMaster_0_M_HADDR(25), 
        ConfigMaster_0_M_HADDR(24) => ConfigMaster_0_M_HADDR(24), 
        ConfigMaster_0_M_HADDR(23) => ConfigMaster_0_M_HADDR(23), 
        ConfigMaster_0_M_HADDR(22) => ConfigMaster_0_M_HADDR(22), 
        ConfigMaster_0_M_HADDR(21) => ConfigMaster_0_M_HADDR(21), 
        ConfigMaster_0_M_HADDR(20) => ConfigMaster_0_M_HADDR(20), 
        ConfigMaster_0_M_HADDR(19) => ConfigMaster_0_M_HADDR(19), 
        ConfigMaster_0_M_HADDR(18) => ConfigMaster_0_M_HADDR(18), 
        ConfigMaster_0_M_HADDR(17) => ConfigMaster_0_M_HADDR(17), 
        ConfigMaster_0_M_HADDR(16) => ConfigMaster_0_M_HADDR(16), 
        ConfigMaster_0_M_HADDR(15) => ConfigMaster_0_M_HADDR(15), 
        ConfigMaster_0_M_HADDR(14) => ConfigMaster_0_M_HADDR(14), 
        ConfigMaster_0_M_HADDR(13) => ConfigMaster_0_M_HADDR(13), 
        ConfigMaster_0_M_HADDR(12) => ConfigMaster_0_M_HADDR(12), 
        ConfigMaster_0_M_HADDR(11) => ConfigMaster_0_M_HADDR(11), 
        ConfigMaster_0_M_HADDR(10) => ConfigMaster_0_M_HADDR(10), 
        ConfigMaster_0_M_HADDR(9) => ConfigMaster_0_M_HADDR(9), 
        ConfigMaster_0_M_HADDR(8) => ConfigMaster_0_M_HADDR(8), 
        ConfigMaster_0_M_HADDR(7) => ConfigMaster_0_M_HADDR(7), 
        ConfigMaster_0_M_HADDR(6) => ConfigMaster_0_M_HADDR(6), 
        ConfigMaster_0_M_HADDR(5) => ConfigMaster_0_M_HADDR(5), 
        ConfigMaster_0_M_HADDR(4) => ConfigMaster_0_M_HADDR(4), 
        ConfigMaster_0_M_HADDR(3) => ConfigMaster_0_M_HADDR(3), 
        ConfigMaster_0_M_HADDR(2) => ConfigMaster_0_M_HADDR(2), 
        ConfigMaster_0_M_HADDR(1) => ConfigMaster_0_M_HADDR(1), 
        ConfigMaster_0_M_HADDR(0) => ConfigMaster_0_M_HADDR(0), 
        ConfigMaster_0_M_HTRANS(1) => ConfigMaster_0_M_HTRANS(1), 
        xhdl1328_i_m_0_1(0) => xhdl1328_i_m_0_1(0), 
        masterDataInProg(0) => masterDataInProg(0), 
        ConfigMaster_0_M_HWDATA(31) => 
        ConfigMaster_0_M_HWDATA(31), ConfigMaster_0_M_HWDATA(30)
         => ConfigMaster_0_M_HWDATA(30), 
        ConfigMaster_0_M_HWDATA(29) => 
        ConfigMaster_0_M_HWDATA(29), ConfigMaster_0_M_HWDATA(28)
         => ConfigMaster_0_M_HWDATA(28), 
        ConfigMaster_0_M_HWDATA(27) => 
        ConfigMaster_0_M_HWDATA(27), ConfigMaster_0_M_HWDATA(26)
         => ConfigMaster_0_M_HWDATA(26), 
        ConfigMaster_0_M_HWDATA(25) => 
        ConfigMaster_0_M_HWDATA(25), ConfigMaster_0_M_HWDATA(24)
         => ConfigMaster_0_M_HWDATA(24), 
        ConfigMaster_0_M_HWDATA(23) => 
        ConfigMaster_0_M_HWDATA(23), ConfigMaster_0_M_HWDATA(22)
         => ConfigMaster_0_M_HWDATA(22), 
        ConfigMaster_0_M_HWDATA(21) => 
        ConfigMaster_0_M_HWDATA(21), ConfigMaster_0_M_HWDATA(20)
         => ConfigMaster_0_M_HWDATA(20), 
        ConfigMaster_0_M_HWDATA(19) => 
        ConfigMaster_0_M_HWDATA(19), ConfigMaster_0_M_HWDATA(18)
         => ConfigMaster_0_M_HWDATA(18), 
        ConfigMaster_0_M_HWDATA(17) => 
        ConfigMaster_0_M_HWDATA(17), ConfigMaster_0_M_HWDATA(16)
         => ConfigMaster_0_M_HWDATA(16), 
        ConfigMaster_0_M_HWDATA(15) => 
        ConfigMaster_0_M_HWDATA(15), ConfigMaster_0_M_HWDATA(14)
         => ConfigMaster_0_M_HWDATA(14), 
        ConfigMaster_0_M_HWDATA(13) => 
        ConfigMaster_0_M_HWDATA(13), ConfigMaster_0_M_HWDATA(12)
         => ConfigMaster_0_M_HWDATA(12), 
        ConfigMaster_0_M_HWDATA(11) => 
        ConfigMaster_0_M_HWDATA(11), ConfigMaster_0_M_HWDATA(10)
         => ConfigMaster_0_M_HWDATA(10), 
        ConfigMaster_0_M_HWDATA(9) => ConfigMaster_0_M_HWDATA(9), 
        ConfigMaster_0_M_HWDATA(8) => ConfigMaster_0_M_HWDATA(8), 
        ConfigMaster_0_M_HWDATA(7) => ConfigMaster_0_M_HWDATA(7), 
        ConfigMaster_0_M_HWDATA(6) => ConfigMaster_0_M_HWDATA(6), 
        ConfigMaster_0_M_HWDATA(5) => ConfigMaster_0_M_HWDATA(5), 
        ConfigMaster_0_M_HWDATA(4) => ConfigMaster_0_M_HWDATA(4), 
        ConfigMaster_0_M_HWDATA(3) => ConfigMaster_0_M_HWDATA(3), 
        ConfigMaster_0_M_HWDATA(2) => ConfigMaster_0_M_HWDATA(2), 
        ConfigMaster_0_M_HWDATA(1) => ConfigMaster_0_M_HWDATA(1), 
        ConfigMaster_0_M_HWDATA(0) => ConfigMaster_0_M_HWDATA(0), 
        CoreAHBLite_1_AHBmslave16_HWDATA(31) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(31), 
        CoreAHBLite_1_AHBmslave16_HWDATA(30) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(30), 
        CoreAHBLite_1_AHBmslave16_HWDATA(29) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(29), 
        CoreAHBLite_1_AHBmslave16_HWDATA(28) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(28), 
        CoreAHBLite_1_AHBmslave16_HWDATA(27) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(27), 
        CoreAHBLite_1_AHBmslave16_HWDATA(26) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(26), 
        CoreAHBLite_1_AHBmslave16_HWDATA(25) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(25), 
        CoreAHBLite_1_AHBmslave16_HWDATA(24) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(24), 
        CoreAHBLite_1_AHBmslave16_HWDATA(23) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(23), 
        CoreAHBLite_1_AHBmslave16_HWDATA(22) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(22), 
        CoreAHBLite_1_AHBmslave16_HWDATA(21) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(21), 
        CoreAHBLite_1_AHBmslave16_HWDATA(20) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(20), 
        CoreAHBLite_1_AHBmslave16_HWDATA(19) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(19), 
        CoreAHBLite_1_AHBmslave16_HWDATA(18) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(18), 
        CoreAHBLite_1_AHBmslave16_HWDATA(17) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(17), 
        CoreAHBLite_1_AHBmslave16_HWDATA(16) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(16), 
        CoreAHBLite_1_AHBmslave16_HWDATA(15) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(15), 
        CoreAHBLite_1_AHBmslave16_HWDATA(14) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(14), 
        CoreAHBLite_1_AHBmslave16_HWDATA(13) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(13), 
        CoreAHBLite_1_AHBmslave16_HWDATA(12) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(12), 
        CoreAHBLite_1_AHBmslave16_HWDATA(11) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(11), 
        CoreAHBLite_1_AHBmslave16_HWDATA(10) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(10), 
        CoreAHBLite_1_AHBmslave16_HWDATA(9) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(9), 
        CoreAHBLite_1_AHBmslave16_HWDATA(8) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(8), 
        CoreAHBLite_1_AHBmslave16_HWDATA(7) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(7), 
        CoreAHBLite_1_AHBmslave16_HWDATA(6) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(6), 
        CoreAHBLite_1_AHBmslave16_HWDATA(5) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(5), 
        CoreAHBLite_1_AHBmslave16_HWDATA(4) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(4), 
        CoreAHBLite_1_AHBmslave16_HWDATA(3) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(3), 
        CoreAHBLite_1_AHBmslave16_HWDATA(2) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(2), 
        CoreAHBLite_1_AHBmslave16_HWDATA(1) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(1), 
        CoreAHBLite_1_AHBmslave16_HWDATA(0) => 
        CoreAHBLite_1_AHBmslave16_HWDATA(0), 
        CoreAHBLite_1_AHBmslave16_HSIZE(1) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(1), 
        CoreAHBLite_1_AHBmslave16_HSIZE(0) => 
        CoreAHBLite_1_AHBmslave16_HSIZE(0), 
        CoreAHBLite_1_AHBmslave16_HADDR(31) => 
        CoreAHBLite_1_AHBmslave16_HADDR(31), 
        CoreAHBLite_1_AHBmslave16_HADDR(30) => 
        CoreAHBLite_1_AHBmslave16_HADDR(30), 
        CoreAHBLite_1_AHBmslave16_HADDR(29) => 
        CoreAHBLite_1_AHBmslave16_HADDR(29), 
        CoreAHBLite_1_AHBmslave16_HADDR(28) => 
        CoreAHBLite_1_AHBmslave16_HADDR(28), 
        CoreAHBLite_1_AHBmslave16_HADDR(27) => 
        CoreAHBLite_1_AHBmslave16_HADDR(27), 
        CoreAHBLite_1_AHBmslave16_HADDR(26) => 
        CoreAHBLite_1_AHBmslave16_HADDR(26), 
        CoreAHBLite_1_AHBmslave16_HADDR(25) => 
        CoreAHBLite_1_AHBmslave16_HADDR(25), 
        CoreAHBLite_1_AHBmslave16_HADDR(24) => 
        CoreAHBLite_1_AHBmslave16_HADDR(24), 
        CoreAHBLite_1_AHBmslave16_HADDR(23) => 
        CoreAHBLite_1_AHBmslave16_HADDR(23), 
        CoreAHBLite_1_AHBmslave16_HADDR(22) => 
        CoreAHBLite_1_AHBmslave16_HADDR(22), 
        CoreAHBLite_1_AHBmslave16_HADDR(21) => 
        CoreAHBLite_1_AHBmslave16_HADDR(21), 
        CoreAHBLite_1_AHBmslave16_HADDR(20) => 
        CoreAHBLite_1_AHBmslave16_HADDR(20), 
        CoreAHBLite_1_AHBmslave16_HADDR(19) => 
        CoreAHBLite_1_AHBmslave16_HADDR(19), 
        CoreAHBLite_1_AHBmslave16_HADDR(18) => 
        CoreAHBLite_1_AHBmslave16_HADDR(18), 
        CoreAHBLite_1_AHBmslave16_HADDR(17) => 
        CoreAHBLite_1_AHBmslave16_HADDR(17), 
        CoreAHBLite_1_AHBmslave16_HADDR(16) => 
        CoreAHBLite_1_AHBmslave16_HADDR(16), 
        CoreAHBLite_1_AHBmslave16_HADDR(15) => 
        CoreAHBLite_1_AHBmslave16_HADDR(15), 
        CoreAHBLite_1_AHBmslave16_HADDR(14) => 
        CoreAHBLite_1_AHBmslave16_HADDR(14), 
        CoreAHBLite_1_AHBmslave16_HADDR(13) => 
        CoreAHBLite_1_AHBmslave16_HADDR(13), 
        CoreAHBLite_1_AHBmslave16_HADDR(12) => 
        CoreAHBLite_1_AHBmslave16_HADDR(12), 
        CoreAHBLite_1_AHBmslave16_HADDR(11) => 
        CoreAHBLite_1_AHBmslave16_HADDR(11), 
        CoreAHBLite_1_AHBmslave16_HADDR(10) => 
        CoreAHBLite_1_AHBmslave16_HADDR(10), 
        CoreAHBLite_1_AHBmslave16_HADDR(9) => 
        CoreAHBLite_1_AHBmslave16_HADDR(9), 
        CoreAHBLite_1_AHBmslave16_HADDR(8) => 
        CoreAHBLite_1_AHBmslave16_HADDR(8), 
        CoreAHBLite_1_AHBmslave16_HADDR(7) => 
        CoreAHBLite_1_AHBmslave16_HADDR(7), 
        CoreAHBLite_1_AHBmslave16_HADDR(6) => 
        CoreAHBLite_1_AHBmslave16_HADDR(6), 
        CoreAHBLite_1_AHBmslave16_HADDR(5) => 
        CoreAHBLite_1_AHBmslave16_HADDR(5), 
        CoreAHBLite_1_AHBmslave16_HADDR(4) => 
        CoreAHBLite_1_AHBmslave16_HADDR(4), 
        CoreAHBLite_1_AHBmslave16_HADDR(3) => 
        CoreAHBLite_1_AHBmslave16_HADDR(3), 
        CoreAHBLite_1_AHBmslave16_HADDR(2) => 
        CoreAHBLite_1_AHBmslave16_HADDR(2), 
        CoreAHBLite_1_AHBmslave16_HADDR(1) => 
        CoreAHBLite_1_AHBmslave16_HADDR(1), 
        CoreAHBLite_1_AHBmslave16_HADDR(0) => 
        CoreAHBLite_1_AHBmslave16_HADDR(0), 
        CoreAHBLite_1_AHBmslave16_HTRANS(1) => 
        CoreAHBLite_1_AHBmslave16_HTRANS(1), HPMS_READY => 
        HPMS_READY, Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, 
        ConfigMaster_0_M_HWRITE => ConfigMaster_0_M_HWRITE, 
        defSlaveSMNextState_m_0_3 => defSlaveSMNextState_m_0_3, 
        un1_state_31_i_i_a2_0_d_1_0_1 => 
        un1_state_31_i_i_a2_0_d_1_0_1, defSlaveSMNextState_m_0_2
         => defSlaveSMNextState_m_0_2, HREADY_i_3 => HREADY_i_3, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, N_98 => N_98, N_25
         => N_25, defSlaveSMNextState_m_0_3_1 => 
        defSlaveSMNextState_m_0_3_1, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, HREADY_i_3_i_0 => HREADY_i_3_i_0, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, 
        CoreAHBLite_1_AHBmslave16_HSELx => 
        CoreAHBLite_1_AHBmslave16_HSELx, 
        CoreAHBLite_1_AHBmslave16_HWRITE => 
        CoreAHBLite_1_AHBmslave16_HWRITE);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreConfigMaster is

    port( ConfigMaster_0_M_HTRANS                 : out   std_logic_vector(1 to 1);
          ConfigMaster_0_M_HWDATA                 : out   std_logic_vector(31 downto 0);
          ConfigMaster_0_M_HSIZE                  : out   std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HRDATA                 : in    std_logic_vector(31 downto 0);
          ConfigMaster_0_M_HADDR                  : out   std_logic_vector(31 downto 0);
          masterDataInProg                        : in    std_logic_vector(0 to 0);
          xhdl1328_i_m_0_1                        : in    std_logic_vector(0 to 0);
          HPMS_READY                              : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          ConfigMaster_0_M_HWRITE                 : out   std_logic;
          HREADY_i_3_i_0                          : in    std_logic;
          defSlaveSMNextState_m_0_3               : in    std_logic;
          defSlaveSMNextState_m_0_2               : in    std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic;
          defSlaveSMNextState_m                   : in    std_logic;
          HREADY_i_3                              : in    std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : in    std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : in    std_logic;
          N_98                                    : in    std_logic;
          N_25                                    : in    std_logic;
          defSlaveSMNextState_m_0_3_1             : in    std_logic
        );

end CoreConfigMaster;

architecture DEF_ARCH of CoreConfigMaster is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \un7_iv_0_a1_0[14]_net_1\, \un7_iv_0_a1_0_i[14]\, 
        VCC_net_1, \un1_state_42_0_0\, \un1_state_46\, GND_net_1, 
        N_727_i_0, N_31, \HWDATA_int_RNO[0]_net_1\, 
        un1_state_38_i_0, \HWDATA_int_RNO[1]_net_1\, 
        \HWDATA_int_RNO[2]_net_1\, \HWDATA_int_RNO[3]_net_1\, 
        \HWDATA_int_RNO[4]_net_1\, \HWDATA_int_RNO[5]_net_1\, 
        \HWDATA_int_RNO[6]_net_1\, \HWDATA_int_RNO[7]_net_1\, 
        \HWDATA_int_RNO[8]_net_1\, \HWDATA_int_RNO[9]_net_1\, 
        N_1897, N_1926, \HWDATA_int_RNO[12]_net_1\, 
        \HWDATA_int_RNO[13]_net_1\, \HWDATA_int_RNO[14]_net_1\, 
        \HWDATA_int_RNO[15]_net_1\, \HWDATA_int_RNO[16]_net_1\, 
        \HWDATA_int_RNO[17]_net_1\, \HWDATA_int_RNO[18]_net_1\, 
        \HWDATA_int_RNO[19]_net_1\, \HWDATA_int_RNO[20]_net_1\, 
        \HWDATA_int_RNO[21]_net_1\, \HWDATA_int_RNO[22]_net_1\, 
        \HWDATA_int_RNO[23]_net_1\, N_2351, 
        \HWDATA_int_RNO[25]_net_1\, \HWDATA_int_RNO[26]_net_1\, 
        \HWDATA_int_RNO[27]_net_1\, \HWDATA_int_RNO[28]_net_1\, 
        \HWDATA_int_RNO[29]_net_1\, N_2525, 
        \HWDATA_int_RNO[31]_net_1\, \haddr_write[0]_net_1\, 
        un46_d_haddr_cry_0_Y, \un1_d_HWRITE_0_sqmuxa_1_0\, 
        \haddr_write[1]_net_1\, un46_d_haddr_cry_1_S, 
        \haddr_write[2]_net_1\, un46_d_haddr_cry_2_S, 
        \haddr_write[3]_net_1\, un46_d_haddr_cry_3_S, 
        \haddr_write[4]_net_1\, un46_d_haddr_cry_4_S, 
        \haddr_write[5]_net_1\, un46_d_haddr_cry_5_S, 
        \haddr_write[6]_net_1\, un46_d_haddr_cry_6_S, 
        \haddr_write[7]_net_1\, un46_d_haddr_cry_7_S, 
        \haddr_write[8]_net_1\, un46_d_haddr_cry_8_S, 
        \haddr_write[9]_net_1\, un46_d_haddr_cry_9_S, 
        \haddr_write[10]_net_1\, un46_d_haddr_cry_10_S, 
        \haddr_write[11]_net_1\, un46_d_haddr_cry_11_S, 
        \haddr_write[12]_net_1\, un46_d_haddr_cry_12_S, 
        \haddr_write[13]_net_1\, un46_d_haddr_cry_13_S, 
        \haddr_write[14]_net_1\, un46_d_haddr_cry_14_S, 
        \haddr_write[15]_net_1\, un46_d_haddr_s_15_S, 
        \haddr_write[16]_net_1\, un46_d_haddr_cry_16_S, 
        \haddr_write[17]_net_1\, un46_d_haddr_cry_17_S, 
        \haddr_write[18]_net_1\, un46_d_haddr_cry_18_S, 
        \haddr_write[19]_net_1\, un46_d_haddr_cry_19_S, 
        \haddr_write[20]_net_1\, un46_d_haddr_cry_20_S, 
        \haddr_write[21]_net_1\, un46_d_haddr_cry_21_S, 
        \haddr_write[22]_net_1\, un46_d_haddr_cry_22_S, 
        \haddr_write[23]_net_1\, un46_d_haddr_cry_23_S, 
        \haddr_write[24]_net_1\, un46_d_haddr_cry_24_S, 
        \haddr_write[25]_net_1\, un46_d_haddr_cry_25_S, 
        \haddr_write[26]_net_1\, un46_d_haddr_cry_26_S, 
        \haddr_write[27]_net_1\, un46_d_haddr_cry_27_S, 
        \haddr_write[28]_net_1\, un46_d_haddr_cry_28_S, 
        \haddr_write[29]_net_1\, un46_d_haddr_cry_29_S, 
        \haddr_write[30]_net_1\, un46_d_haddr_cry_30_S, 
        \haddr_write[31]_net_1\, un46_d_haddr_s_31_S, 
        \ins2[0]_net_1\, \d_ins2[0]_net_1\, N_654, 
        \ins2[1]_net_1\, \d_ins2[1]_net_1\, \ins2[2]_net_1\, 
        \d_ins2[2]_net_1\, \ins2[3]_net_1\, \d_ins2[3]_net_1\, 
        \ins2[4]_net_1\, \d_ins2[4]_net_1\, \ins2[5]_net_1\, 
        \d_ins2[5]_net_1\, \ins2[6]_net_1\, \d_ins2[6]_net_1\, 
        \ins2[7]_net_1\, \d_ins2[7]_net_1\, \ins2[8]_net_1\, 
        \d_ins2[8]_net_1\, \ins2[9]_net_1\, \d_ins2[9]_net_1\, 
        \ins2[10]_net_1\, \d_ins2[10]_net_1\, \ins2[11]_net_1\, 
        \d_ins2[11]_net_1\, \ins2[12]_net_1\, \d_ins2[12]_net_1\, 
        \ins2[13]_net_1\, \d_ins2[13]_net_1\, \ins2[14]_net_1\, 
        \d_ins2[14]_net_1\, \ins2[15]_net_1\, \d_ins2[15]_net_1\, 
        \ins2[16]_net_1\, \d_ins2[16]_net_1\, \ins2[17]_net_1\, 
        \d_ins2[17]_net_1\, \ins2[18]_net_1\, \d_ins2[18]_net_1\, 
        \ins2[19]_net_1\, \d_ins2[19]_net_1\, \ins2[20]_net_1\, 
        \d_ins2[20]_net_1\, \ins2[21]_net_1\, \d_ins2[21]_net_1\, 
        \ins2[22]_net_1\, \d_ins2[22]_net_1\, \ins2[23]_net_1\, 
        \d_ins2[23]_net_1\, \ins2[24]_net_1\, \d_ins2[24]_net_1\, 
        \ins2[25]_net_1\, \d_ins2[25]_net_1\, \ins2[26]_net_1\, 
        \d_ins2[26]_net_1\, \ins2[27]_net_1\, \d_ins2[27]_net_1\, 
        \ins2[28]_net_1\, \d_ins2[28]_net_1\, \ins2[29]_net_1\, 
        \d_ins2[29]_net_1\, \ins2[30]_net_1\, \d_ins2[30]_net_1\, 
        \ins2[31]_net_1\, \d_ins2[31]_net_1\, N_415, 
        \un1_state_34_0_0\, \acc[0]_net_1\, \d_acc[0]\, 
        \un1_state_25_0_0\, \acc[1]_net_1\, \d_acc[1]_net_1\, 
        \acc[2]_net_1\, \d_acc[2]_net_1\, \acc[3]_net_1\, 
        \d_acc[3]\, \acc[4]_net_1\, \d_acc[4]\, \acc[5]_net_1\, 
        \d_acc[5]\, \acc[6]_net_1\, \d_acc[6]_net_1\, 
        \acc[7]_net_1\, \d_acc[7]\, \acc[8]_net_1\, 
        \d_acc[8]_net_1\, \acc[9]_net_1\, \d_acc[9]_net_1\, 
        \acc[10]_net_1\, \d_acc[10]\, \acc[11]_net_1\, 
        \d_acc[11]_net_1\, \acc[12]_net_1\, \d_acc[12]_net_1\, 
        \acc[13]_net_1\, \d_acc[13]\, \acc[14]_net_1\, 
        \d_acc[14]_net_1\, \acc[15]_net_1\, \d_acc[15]_net_1\, 
        \acc[16]_net_1\, \d_acc[16]\, \acc[17]_net_1\, 
        \d_acc[17]_net_1\, \acc[18]_net_1\, \d_acc[18]\, 
        \acc[19]_net_1\, \d_acc[19]_net_1\, \acc[20]_net_1\, 
        \d_acc[20]_net_1\, \acc[21]_net_1\, \d_acc[21]\, 
        \acc[22]_net_1\, \d_acc[22]_net_1\, \acc[23]_net_1\, 
        \d_acc[23]_net_1\, \acc[24]_net_1\, \d_acc[24]\, 
        \acc[25]_net_1\, \d_acc[25]_net_1\, \acc[26]_net_1\, 
        \d_acc[26]_net_1\, \acc[27]_net_1\, \d_acc[27]_net_1\, 
        \acc[28]_net_1\, \d_acc[28]\, \acc[29]_net_1\, 
        \d_acc[29]_net_1\, \acc[30]_net_1\, \d_acc[30]\, 
        \acc[31]_net_1\, \d_acc[31]_net_1\, \busy\, d_busy, 
        \state[2]_net_1\, \rdata[0]_net_1\, N_725_i_0, 
        \rdata[1]_net_1\, \rdata[2]_net_1\, \rdata[3]_net_1\, 
        \rdata[4]_net_1\, \rdata[5]_net_1\, \rdata[6]_net_1\, 
        \rdata[7]_net_1\, \rdata[8]_net_1\, \rdata[9]_net_1\, 
        \rdata[10]_net_1\, \rdata[11]_net_1\, \rdata[12]_net_1\, 
        \rdata[13]_net_1\, \rdata[14]_net_1\, \rdata[15]_net_1\, 
        \rdata[16]_net_1\, \rdata[17]_net_1\, \rdata[18]_net_1\, 
        \rdata[19]_net_1\, \rdata[20]_net_1\, \rdata[21]_net_1\, 
        \rdata[22]_net_1\, \rdata[23]_net_1\, \rdata[24]_net_1\, 
        \rdata[25]_net_1\, \rdata[26]_net_1\, \rdata[27]_net_1\, 
        \rdata[28]_net_1\, \rdata[29]_net_1\, \rdata[30]_net_1\, 
        \rdata[31]_net_1\, \mask[0]_net_1\, N_167, 
        \mask[1]_net_1\, \mask[2]_net_1\, \mask[3]_net_1\, 
        \mask[4]_net_1\, \mask[5]_net_1\, \mask[6]_net_1\, 
        \mask[7]_net_1\, \mask[8]_net_1\, \mask[9]_net_1\, 
        \mask[10]_net_1\, \mask[11]_net_1\, \mask[12]_net_1\, 
        \mask[13]_net_1\, \mask[14]_net_1\, \mask[15]_net_1\, 
        \mask[16]_net_1\, \mask[17]_net_1\, \mask[18]_net_1\, 
        \mask[19]_net_1\, \mask[20]_net_1\, \mask[21]_net_1\, 
        \mask[22]_net_1\, \mask[23]_net_1\, \mask[24]_net_1\, 
        \mask[25]_net_1\, \mask[26]_net_1\, \mask[27]_net_1\, 
        \mask[28]_net_1\, \mask[29]_net_1\, \mask[30]_net_1\, 
        \mask[31]_net_1\, \ins1[0]_net_1\, N_700_i_0, 
        \ins1[1]_net_1\, \ins1[2]_net_1\, \ins1[3]_net_1\, 
        \ins1[4]_net_1\, \ins1[5]_net_1\, \ins1[6]_net_1\, 
        \ins1[7]_net_1\, \ins1[8]_net_1\, \ins1[9]_net_1\, 
        \ins1[10]_net_1\, \ins1[11]_net_1\, \ins1[12]_net_1\, 
        \ins1[13]_net_1\, \ins1[14]_net_1\, \ins1[15]_net_1\, 
        \ins1[16]_net_1\, \ins1[17]_net_1\, \ins1[18]_net_1\, 
        \ins1[19]_net_1\, \ins1[20]_net_1\, \ins1[21]_net_1\, 
        \ins1[22]_net_1\, \ins1[23]_net_1\, \ins1[24]_net_1\, 
        \ins1[25]_net_1\, \ins1[26]_net_1\, \ins1[27]_net_1\, 
        \ins1[28]_net_1\, \ins1[29]_net_1\, \ins1[30]_net_1\, 
        \ins1[31]_net_1\, \expected[0]_net_1\, N_702_i_0, 
        \expected[1]_net_1\, \expected[2]_net_1\, 
        \expected[3]_net_1\, \expected[4]_net_1\, 
        \expected[5]_net_1\, \expected[6]_net_1\, 
        \expected[7]_net_1\, \expected[8]_net_1\, 
        \expected[9]_net_1\, \expected[10]_net_1\, 
        \expected[11]_net_1\, \expected[12]_net_1\, 
        \expected[13]_net_1\, \expected[14]_net_1\, 
        \expected[15]_net_1\, \expected[16]_net_1\, 
        \expected[17]_net_1\, \expected[18]_net_1\, 
        \expected[19]_net_1\, \expected[20]_net_1\, 
        \expected[21]_net_1\, \expected[22]_net_1\, 
        \expected[23]_net_1\, \expected[24]_net_1\, 
        \expected[25]_net_1\, \expected[26]_net_1\, 
        \expected[27]_net_1\, \expected[28]_net_1\, 
        \expected[29]_net_1\, \expected[30]_net_1\, 
        \expected[31]_net_1\, \envm_soft_reset[0]_net_1\, 
        N_696_i_0, \envm_soft_reset[1]_net_1\, 
        \envm_busy[0]_net_1\, N_14_i_0, \envm_busy[1]_net_1\, 
        \pause_count[2]_net_1\, N_4807_i_0, pause_counte, 
        \pause_count[3]_net_1\, N_4808_i_0, 
        \pause_count[4]_net_1\, N_4809_i_0, 
        \pause_count[0]_net_1\, N_4316_i_0, 
        \pause_count[1]_net_1\, N_37_i_0, \bytecount[13]_net_1\, 
        N_52_i_0, \bytecount[14]_net_1\, N_55_i_0, 
        \bytecount[15]_net_1\, \d_bytecount[15]_net_1\, 
        \count[0]_net_1\, N_4888_i_0, \count[1]_net_1\, 
        \d_count[1]\, \bytecount[0]_net_1\, N_28_i_0, 
        \bytecount[1]_net_1\, \d_bytecount[1]_net_1\, 
        \bytecount[2]_net_1\, N_32_i_0, \bytecount[3]_net_1\, 
        \d_bytecount[3]_net_1\, \bytecount[4]_net_1\, N_34_i_0, 
        \bytecount[5]_net_1\, N_36_i_0, \bytecount[6]_net_1\, 
        N_38_i_0, \bytecount[7]_net_1\, N_40_i_0, 
        \bytecount[8]_net_1\, N_42_i_0, \bytecount[9]_net_1\, 
        N_44_i_0, \bytecount[10]_net_1\, N_46_i_0, 
        \bytecount[11]_net_1\, N_48_i_0, \bytecount[12]_net_1\, 
        N_50_i_0, \haddr_fetch[17]_net_1\, N_4403_i_0, 
        \un1_d_haddr_fetch_2_sqmuxa\, \haddr_fetch[18]_net_1\, 
        \haddr_fetch_RNO[18]_net_1\, \haddr_fetch[19]_net_1\, 
        N_4367_i_0, \haddr_fetch[20]_net_1\, N_4560_i_0, 
        \haddr_fetch[21]_net_1\, N_62, \haddr_fetch[22]_net_1\, 
        N_4722_i_0, \haddr_fetch[23]_net_1\, N_3216_i_0, 
        \haddr_fetch[24]_net_1\, \haddr_fetch_RNO[24]_net_1\, 
        \haddr_fetch[25]_net_1\, N_3162_i_0, 
        \haddr_fetch[26]_net_1\, N_21_i_0, 
        \haddr_fetch[27]_net_1\, N_4407_i_0, 
        \haddr_fetch[28]_net_1\, N_19_i_0, 
        \haddr_fetch[29]_net_1\, N_18_i_0, 
        \haddr_fetch[30]_net_1\, N_17_i_0, 
        \haddr_fetch[31]_net_1\, N_4366_i_0, 
        \haddr_fetch[2]_net_1\, N_64_i, \haddr_fetch[3]_net_1\, 
        N_53_i_0, \haddr_fetch[4]_net_1\, N_2921_i_0, 
        \haddr_fetch[5]_net_1\, \haddr_fetch_RNO[5]_net_1\, 
        \haddr_fetch[6]_net_1\, N_4720_i_0, 
        \haddr_fetch[7]_net_1\, \haddr_fetch_RNO[7]_net_1\, 
        \haddr_fetch[8]_net_1\, N_4365_i_0, 
        \haddr_fetch[9]_net_1\, N_4418_i_0, 
        \haddr_fetch[10]_net_1\, N_4364_i_0, 
        \haddr_fetch[11]_net_1\, N_119_i_0, 
        \haddr_fetch[12]_net_1\, N_4402_i_0, 
        \haddr_fetch[13]_net_1\, \haddr_fetch_RNO[13]_net_1\, 
        \haddr_fetch[14]_net_1\, N_2651_i_0, 
        \haddr_fetch[15]_net_1\, N_4342_i_0, 
        \haddr_fetch[16]_net_1\, N_4719_i_0, 
        \haddr_fetch[0]_net_1\, \ConfigMaster_0_M_HADDR[0]\, 
        \haddr_fetch[1]_net_1\, \ConfigMaster_0_M_HADDR[1]\, 
        \ConfigMaster_0_M_HADDR[24]\, \d_HADDR[24]\, 
        un1_state_44_i_0, \ConfigMaster_0_M_HADDR[25]\, 
        \d_HADDR[25]\, \ConfigMaster_0_M_HADDR[26]\, 
        \d_HADDR[26]\, \ConfigMaster_0_M_HADDR[27]\, 
        \d_HADDR[27]\, \ConfigMaster_0_M_HADDR[28]\, 
        \d_HADDR[28]\, \ConfigMaster_0_M_HADDR[29]\, 
        \d_HADDR[29]\, \ConfigMaster_0_M_HADDR[30]\, 
        \d_HADDR_0_iv_i_0[30]\, \ConfigMaster_0_M_HADDR[31]\, 
        \d_HADDR[31]\, \ConfigMaster_0_M_HADDR[9]\, \d_HADDR[9]\, 
        \ConfigMaster_0_M_HADDR[10]\, \d_HADDR[10]\, 
        \ConfigMaster_0_M_HADDR[11]\, \d_HADDR[11]\, 
        \ConfigMaster_0_M_HADDR[12]\, \d_HADDR[12]\, 
        \ConfigMaster_0_M_HADDR[13]\, \d_HADDR[13]\, 
        \ConfigMaster_0_M_HADDR[14]\, \d_HADDR[14]\, 
        \ConfigMaster_0_M_HADDR[15]\, \d_HADDR_0_iv_i_0[15]\, 
        \ConfigMaster_0_M_HADDR[16]\, \d_HADDR_0_iv_i_0[16]\, 
        \ConfigMaster_0_M_HADDR[17]\, \d_HADDR_0_iv_i_0[17]\, 
        \ConfigMaster_0_M_HADDR[18]\, \d_HADDR[18]\, 
        \ConfigMaster_0_M_HADDR[19]\, \d_HADDR[19]\, 
        \ConfigMaster_0_M_HADDR[20]\, \d_HADDR[20]\, 
        \ConfigMaster_0_M_HADDR[21]\, \d_HADDR[21]\, 
        \ConfigMaster_0_M_HADDR[22]\, \d_HADDR[22]\, 
        \ConfigMaster_0_M_HADDR[23]\, \d_HADDR[23]\, \d_HADDR[0]\, 
        \d_HADDR[1]\, \ConfigMaster_0_M_HADDR[2]\, \d_HADDR[2]\, 
        \ConfigMaster_0_M_HADDR[3]\, \d_HADDR_0_iv_i_0[3]\, 
        \ConfigMaster_0_M_HADDR[4]\, \d_HADDR[4]\, 
        \ConfigMaster_0_M_HADDR[5]\, \d_HADDR[5]\, 
        \ConfigMaster_0_M_HADDR[6]\, \d_HADDR_0_iv_i_0[6]\, 
        \ConfigMaster_0_M_HADDR[7]\, \d_HADDR[7]\, 
        \ConfigMaster_0_M_HADDR[8]\, \d_HADDR[8]\, 
        \state[4]_net_1\, \state_ns[24]\, \state[3]_net_1\, 
        \state[1]_net_1\, \state[0]_net_1\, \state_ns[28]\, 
        \state[19]_net_1\, \state_ns[9]\, \state[18]_net_1\, 
        \state[17]_net_1\, \state_ns[11]\, \state[16]_net_1\, 
        N_480, \state[15]_net_1\, \state_ns[13]\, 
        \state[14]_net_1\, N_16_i_0, \state[13]_net_1\, 
        \state[12]_net_1\, \state_ns[16]_net_1\, 
        \state[11]_net_1\, \state_ns[17]\, \state[10]_net_1\, 
        \state[9]_net_1\, \state[8]_net_1\, \state_ns[20]\, 
        \state[7]_net_1\, N_20_i_0, \state[6]_net_1\, 
        \state_ns[22]\, \state[5]_net_1\, \state[28]_net_1\, 
        \state_ns[0]\, \state[27]_net_1\, N_741_i_0, 
        \state[26]_net_1\, \state_ns[2]\, \state[25]_net_1\, 
        N_70_i_0, \state[24]_net_1\, N_12_i_0, \state[23]_net_1\, 
        \state_ns[5]\, \state[22]_net_1\, N_170, 
        \state[21]_net_1\, \state_ns[7]\, \state[20]_net_1\, 
        \state_ns[8]\, \HADDR_int_fast[0]_net_1\, 
        \d_HADDR_fast[0]\, \state_fast[21]_net_1\, 
        \state_ns_fast[7]\, \state_21_rep1\, \state_ns_rep1[7]\, 
        un13_d_haddr_1_cry_27_1_FCO, un13_d_haddr_1_cry_27_3_FCO, 
        un13_d_haddr_1_cry_27_5_FCO, \un13_d_haddr_1_cry_13\, 
        un13_d_haddr_1_cry_13_S, \un13_d_haddr_1_cry_14\, 
        un13_d_haddr_1_cry_14_S, \un13_d_haddr_1_cry_15\, 
        un13_d_haddr_1_cry_15_S, \un13_d_haddr_1_cry_16\, 
        un13_d_haddr_1_cry_16_S, \un13_d_haddr_1_cry_17\, 
        un13_d_haddr_1_cry_17_S, \un13_d_haddr_1_cry_18\, 
        un13_d_haddr_1_cry_18_S, \un13_d_haddr_1_cry_19\, 
        un13_d_haddr_1_cry_19_S, \un13_d_haddr_1_cry_20\, 
        un13_d_haddr_1_cry_20_S, \un13_d_haddr_1_cry_21\, 
        un13_d_haddr_1_cry_21_S, \un13_d_haddr_1_cry_22\, 
        un13_d_haddr_1_cry_22_S, \un13_d_haddr_1_cry_23\, 
        un13_d_haddr_1_cry_23_S, \un13_d_haddr_1_cry_24\, 
        un13_d_haddr_1_cry_24_S, \un13_d_haddr_1_cry_25\, 
        un13_d_haddr_1_cry_25_S, \un13_d_haddr_1_cry_26\, 
        un13_d_haddr_1_cry_26_S, \un13_d_haddr_1_cry_27\, 
        un13_d_haddr_1_cry_27_S, un13_d_haddr_1_s_29_S, 
        \un13_d_haddr_1_cry_28\, un13_d_haddr_1_cry_28_S, 
        un46_d_haddr_cry_0_0_FCO, un46_d_haddr_cry_1_0_FCO, 
        un46_d_haddr_cry_2_0_FCO, un46_d_haddr_cry_3_0_FCO, 
        un46_d_haddr_cry_30_1_FCO, un46_d_haddr_cry_30_3_FCO, 
        un46_d_haddr_cry_30_5_FCO, \un46_d_haddr_cry_16\, 
        \un46_d_haddr_cry_17\, \un46_d_haddr_cry_18\, 
        \un46_d_haddr_cry_19\, \un46_d_haddr_cry_20\, 
        \un46_d_haddr_cry_21\, \un46_d_haddr_cry_22\, 
        \un46_d_haddr_cry_23\, \un46_d_haddr_cry_24\, 
        \un46_d_haddr_cry_25\, \un46_d_haddr_cry_26\, 
        \un46_d_haddr_cry_27\, \un46_d_haddr_cry_28\, 
        \un46_d_haddr_cry_29\, \un46_d_haddr_cry_30\, 
        d_bytecount_i_m2_cry_0, \ins1_RNIE4ISO_Y[0]\, N_78, N_166, 
        d_bytecount_i_m2_cry_1, N_1102, \un7_iv[14]_net_1\, 
        d_bytecount_i_m2_cry_2, N_104, N_164, 
        d_bytecount_i_m2_cry_3, N_1104, d_bytecount_i_m2_cry_4, 
        N_105, d_bytecount_i_m2_cry_5, N_106, 
        d_bytecount_i_m2_cry_6, N_4336, d_bytecount_i_m2_cry_7, 
        N_108, d_bytecount_i_m2_cry_8, N_4337, 
        d_bytecount_i_m2_cry_9, N_4338, d_bytecount_i_m2_cry_10, 
        N_4339, d_bytecount_i_m2_cry_11, N_4340, 
        d_bytecount_i_m2_cry_12, N_114, d_bytecount_i_m2_cry_13, 
        N_4341, N_1116, d_bytecount_i_m2_cry_14, N_116, 
        \un46_d_haddr_cry_0\, \un46_d_haddr_cry_1\, 
        \un46_d_haddr_cry_2\, \un46_d_haddr_cry_3\, 
        \un46_d_haddr_cry_4\, \un46_d_haddr_cry_5\, 
        \un46_d_haddr_cry_6\, \un46_d_haddr_cry_7\, 
        \un46_d_haddr_cry_8\, \un46_d_haddr_cry_9\, 
        \un46_d_haddr_cry_10\, \un46_d_haddr_cry_11\, 
        \un46_d_haddr_cry_12\, \un46_d_haddr_cry_13\, 
        \un46_d_haddr_cry_14\, \un1_rdata_0_data_tmp[0]\, N_83_i, 
        \un1_rdata_0_data_tmp[1]\, N_347_i, 
        \un1_rdata_0_data_tmp[2]\, un1_rdata_0_N_12, 
        \un1_rdata_0_data_tmp[3]\, un1_rdata_0_N_57, 
        \un1_rdata_0_data_tmp[4]\, un1_rdata_0_N_37, 
        \un1_rdata_0_data_tmp[5]\, N_351_i, 
        \un1_rdata_0_data_tmp[6]\, N_343_i, 
        \un1_rdata_0_data_tmp[7]\, N_339_i, 
        \un1_rdata_0_data_tmp[8]\, N_323_i, 
        \un1_rdata_0_data_tmp[9]\, N_335_i, 
        \un1_rdata_0_data_tmp[10]\, un1_rdata_0_N_53, 
        \un1_rdata_0_data_tmp[11]\, N_359_i, 
        \un1_rdata_0_data_tmp[12]\, N_327_i, 
        \un1_rdata_0_data_tmp[13]\, N_331_i, 
        \un1_rdata_0_data_tmp[14]\, N_355_i, d_state61_li, 
        un1_rdata_0_N_22, un13_d_haddr_1_s_1_172_FCO, 
        \un13_d_haddr_1_cry_1\, un13_d_haddr_1_cry_1_S, 
        \un13_d_haddr_1_cry_2\, un13_d_haddr_1_cry_2_S, 
        \un13_d_haddr_1_cry_3\, un13_d_haddr_1_cry_3_S, 
        \un13_d_haddr_1_cry_4\, un13_d_haddr_1_cry_4_S, 
        \un13_d_haddr_1_cry_5\, un13_d_haddr_1_cry_5_S, 
        \un13_d_haddr_1_cry_6\, un13_d_haddr_1_cry_6_S, 
        \un13_d_haddr_1_cry_7\, un13_d_haddr_1_cry_7_S, 
        \un13_d_haddr_1_cry_8\, un13_d_haddr_1_cry_8_S, 
        \un13_d_haddr_1_cry_9\, un13_d_haddr_1_cry_9_S, 
        \un13_d_haddr_1_cry_10\, un13_d_haddr_1_cry_10_S, 
        un13_d_haddr_1_s_12_S, \un13_d_haddr_1_cry_11\, 
        un13_d_haddr_1_cry_11_S, \un1_state_44_0_6\, 
        \un1_state_44_0_4\, \un1_state_44_0_8\, 
        \un1_state_44_0_9\, un1_state_31_i_i_a2_0_d_1_sx_0, 
        un1_state_31_i_i_a2_0_d_1_0_sx, N_290, 
        un1_state_31_i_i_o2_0, d_state_1_sqmuxa_1_i_0, N_109_i, 
        N_101, \un1_state_30_0_0\, \d_HADDR_0_iv_1_1[31]_net_1\, 
        N_4814, \d_HADDR_0_iv_1_0[31]_net_1\, N_247, 
        un1_d_HWRITE_0_sqmuxa_2, \d_HADDR_0_iv_0_2[0]_net_1\, 
        \d_HADDR_0_iv_0_2[30]_net_1\, \d_HADDR_0_iv_i_1[30]\, 
        \d_HADDR_0_iv_0_0[30]_net_1\, 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, \un13_d_haddr_1_i_m[15]\, 
        \d_HADDR_0_iv_i_1[15]\, \d_HADDR_0_iv_1[15]_net_1\, 
        \d_HADDR_0_iv_0_2[3]_net_1\, \d_HADDR_0_iv_i_1[3]\, 
        \d_HADDR_0_iv_0_0[3]_net_1\, \d_HADDR_0_iv_2[6]_net_1\, 
        \d_HADDR_0_iv_i_1[6]\, \d_HADDR_0_iv_0[6]_net_1\, 
        \un13_d_haddr_1_m[29]\, \d_HADDR_0_iv_1_0[29]_net_1\, 
        \d_HADDR_0_iv_1[29]_net_1\, \un13_d_haddr_1_m[27]\, 
        \d_HADDR_0_iv_1_0[27]_net_1\, \d_HADDR_0_iv_1[27]_net_1\, 
        \d_HADDR_0_iv_0_2[13]_net_1\, 
        \d_HADDR_0_iv_0_1[13]_net_1\, 
        \d_HADDR_0_iv_0_0[13]_net_1\, \d_HADDR_0_iv_0_1[7]_net_1\, 
        \d_HADDR_0_iv_0_1_0[7]_net_1\, N_4592, 
        \d_HADDR_0_iv_2[14]_net_1\, \d_HADDR_0_iv_1[14]_net_1\, 
        \d_HADDR_0_iv_0[14]_net_1\, \un13_d_haddr_1_m[1]\, 
        \d_HADDR_0_iv_1_0[1]_net_1\, \d_HADDR_0_iv_1[1]_net_1\, 
        \d_HADDR_0_iv_1[31]_net_1\, \d_HADDR_0_iv_2[8]_net_1\, 
        \d_HADDR_0_iv_1[8]_net_1\, \d_HADDR_0_iv_0[8]_net_1\, 
        \un13_d_haddr_1_m[22]\, \d_HADDR_0_iv_1_0[22]_net_1\, 
        \d_HADDR_0_iv_1[22]_net_1\, \d_HADDR_0_iv_2[4]_net_1\, 
        \d_HADDR_0_iv_1[4]_net_1\, \d_HADDR_0_iv_0[4]_net_1\, 
        \d_HADDR_0_iv_2[11]_net_1\, \d_HADDR_0_iv_1[11]_net_1\, 
        \d_HADDR_0_iv_0[11]_net_1\, 
        \d_HADDR_0_iv_0_0_0[24]_net_1\, 
        \d_HADDR_0_iv_0_0_1[24]_net_1\, N_481, N_252, d_N_3_mux_0, 
        N_294, \d_count_0_o2_0_1_2[1]\, N_445, N_319, N_259, 
        N_375, d_m2_e_2_2, N_4901, N_4902, 
        \un1_d_HWRITE_1_sqmuxa_2_i_o2_1\, N_251, 
        un1_d_HWRITE_1_sqmuxa_2_i_o3_1_2, N_86, 
        \state_ns_i_0_a2_3_0_1[1]_net_1\, N_93_i, N_74, N_917, 
        N_156, N_117, \state_ns_i_a2_10_i_2[1]_net_1\, 
        \d_count_i_a2_2_1_0[0]\, \d_count_i_a2_2_1[0]\, N_452, 
        N_542_2, \d_count_0_a3_8_0[1]\, d_m2_e_1, d_m2_e_2_0_1, 
        d_m2_e_2_0, \un7_iv_1[14]_net_1\, 
        un1_state_31_i_i_a2_0_d_0_0_0, 
        \un1_state_31_i_i_a2_0_d_0_0_1\, d_HWDATA_0_iv_0_1604_5_0, 
        N_4778, d_HWDATA_0_iv_0_1604_1_0, N_680_2, N_4777_1, 
        N_403, d_HWDATA_0_iv_1640_1, N_2061, N_276, 
        d_HWDATA_0_iv_1640_2, N_2573_1, N_272, 
        d_HWDATA_0_iv_14_1028_0_a2_i_1, N_317, N_178, N_249, 
        d_HWDATA_0_iv_1640_2_1, N_2579, d_HWDATA_0_iv_1640_a8_3_0, 
        N_2066, \state_ns_i_a2_13_0_a3_5_0[1]_net_1\, 
        \un1_state_39_3\, \state_ns_i_a2_13_0_a3_5[1]_net_1\, 
        d_HWDATA_0_iv_8_1298_1_o2_i_m2_ns_1, N_390, 
        \d_count_0_a2_1_2_1[1]\, N_541, \d_count_0_a2_1_d[1]\, 
        d_HWDATA_0_iv_11_1163_0_0, N_288, N_283, 
        \d_count_0_o2_0[1]\, N_281, 
        \d_HADDR_0_iv_0_0_a3_0_0[24]_net_1\, 
        \d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0\, 
        d_HWDATA_0_iv_5_1424_a8_0_0, \un9_opcode_0_a2_0\, 
        \d_acc_1_a2_0_0[5]\, \d_HTRANS_0_sqmuxa_4_1_1_o3_1\, 
        \un46_d_haddr_axb_0\, un9_hready_2, N_138, N_475, N_485, 
        N_585, N_263, N_266, N_274, N_4812, N_661, N_4711, N_4539, 
        N_4541, N_200, N_789, N_4912, N_3400, N_125, N_2570, 
        N_388, \state_m3_i_2\, \state_ns_0_a3_2_3[8]_net_1\, 
        \state_ns_0_a3_2_2[8]_net_1\, 
        \un1_d_HWRITE_1_sqmuxa_2_i_o3_0\, 
        \state_ns_i_a2_10_i_1[1]_net_1\, \d_count_0_a3_3_0[1]\, 
        d_m1_e_1_1, \un12_size_2_0_5\, \un12_size_2_0_4\, 
        \un1_state_39_1_0_a3_0_1\, N_80, N_837, N_369, N_4472, 
        N_4811, N_66_i, \state_ns_0_0[8]_net_1\, 
        \un1_state_42_0_0_1\, d_HWDATA_0_iv_3_1496_0_0, 
        d_HWDATA_0_iv_4_1460_5_0, \d_count_0_a3_13_0[1]\, 
        d_HWDATA_0_iv_9_1253_1_0, d_HWDATA_0_iv_25_605_7_0, 
        d_HWDATA_0_iv_5_1424_0, d_HWDATA_0_iv_15_992_0, 
        \d_acc_1_0[0]_net_1\, \d_acc_1_0_0[24]_net_1\, 
        \d_acc_1_0[16]_net_1\, \d_acc_1_0[21]_net_1\, 
        \d_acc_1_0[28]_net_1\, \d_acc_1_0[30]_net_1\, 
        \d_acc_1_0[18]_net_1\, \d_acc_1_0[4]_net_1\, 
        \d_acc_1_0[10]_net_1\, \d_acc_1_0_0[7]_net_1\, 
        \d_acc_1_0[3]_net_1\, \d_acc_1_0[5]_net_1\, 
        \d_acc_1_0[13]_net_1\, \un1_d_HWRITE_0_sqmuxa_0_1\, 
        N_4741, N_465, N_4885, \d_HWRITE_0_sqmuxa_1_0_a3_1\, 
        \d_HTRANS_0_sqmuxa_4_1\, \d_count_0_a2_2_0[1]\, N_133, 
        N_136, N_137, N_591, \un1_state_39_1\, 
        \state_ns_0_a3_2[8]_net_1\, 
        un1_d_HWRITE_1_sqmuxa_2_i_o3_1_0, \d_count_i_a2_1_0[0]\, 
        d_HWDATA_0_iv_9_1253_1_1, d_HWDATA_0_iv_25_605_7_1, 
        d_HWDATA_0_iv_5_1424_1, d_HWDATA_0_iv_25_605_7_1_0, 
        d_HWDATA_0_iv_7_1343_o2_0_0, \un1_d_HWRITE_0_sqmuxa_0_2\, 
        d_HWDATA_0_iv_20_812_o3_0_0, 
        d_HWDATA_0_iv_14_1028_2_a2_i_1, N_2063, N_4917, 
        \d_count_0_0_tz[1]\, N_4525, N_255, N_258, N_4916, N_656, 
        N_4625, N_4653, N_4879, N_512_1, N_4687, N_97, N_198, 
        N_4813, \un1_state_44_0_10\, \d_count_0_o3_3_0[1]\, 
        \un1_d_HWRITE_0_sqmuxa_5_i_a3_1_0\, 
        \d_haddr_fetch_2_sqmuxa_0\, d_HWDATA_0_iv_15_992_2, 
        d_HWDATA_0_iv_8_1298_1_0, d_HWDATA_0_iv_25_605_7_1_1, 
        d_HWDATA_0_iv_8_1298_1_o2_i_1, N_2400, N_2060, N_4889, 
        N_4431, N_257, N_47, N_592, N_601, N_674, N_262, N_291, 
        N_4890, N_4855, N_191, N_543, \state_m3_i_4\, 
        \state_m2_e_0\, d_HWDATA_0_iv_3_1496_0_2, 
        \state_ns_0_a2_0_1[5]_net_1\, 
        \un1_d_HWRITE_1_sqmuxa_2_i_a2_0_0\, 
        \un1_d_HWRITE_0_sqmuxa_1_0_a3_i_1\, un1_m3_e_1, 
        d_HWDATA_0_iv_15_992_4, d_HWDATA_0_iv_30_380_1_0, 
        d_HWDATA_0_iv_14_1028_3_1, 
        \state_ns_i_a2_13_0_a3_8[1]_net_1\, 
        d_HWDATA_0_iv_24_650_7_0, N_2399, N_4891, N_4577, N_579, 
        N_404, un28_opcode, N_402, N_379, N_2380_3, N_587, N_655, 
        N_270, N_271, N_277, N_301, N_254, d_HWRITE_0_sqmuxa_2, 
        N_1146, N_1148, N_1151, N_1157, N_1145, N_1149, N_1154, 
        N_1162, N_1163, N_1168, N_1138, N_1139, N_1152, N_1143, 
        N_1156, N_1159, N_1164, \un1_d_state_1_sqmuxa_1[0]\, 
        N_1160, N_1166, \d_count_i_0[0]\, 
        d_HWDATA_0_iv_10_1208_0_1, d_HWDATA_0_iv_13_1073_0_1, 
        d_HWDATA_0_iv_7_1343_1_0, d_HWDATA_0_iv_12_1118_0_0, 
        d_HWDATA_0_iv_4_1460_5_2, \un1_hready_2_0_0\, 
        d_HWDATA_0_iv_30_380_1_2, N_2246_1, 
        \un1_d_HWRITE_0_sqmuxa\, N_600, N_264, N_278, 
        \d_count_i_1[0]\, un1_d_HWRITE_0_sqmuxa_5_i_a3_0, 
        d_HWDATA_0_iv_26_560_0_0, d_HWDATA_0_iv_27_515_0_0, 
        d_HWDATA_0_iv_23_695_0_0, d_HWDATA_0_iv_28_470_3_0, 
        d_HWDATA_0_iv_29_425_0_0, d_HWDATA_0_iv_18_884_6_0, 
        d_HWDATA_0_iv_22_740_6_0, d_HWDATA_0_iv_19_848_6_0, 
        d_HWDATA_0_iv_20_812_0_0, d_HWDATA_0_iv_16_956_0_0, 
        d_HWDATA_0_iv_21_776_6_0, d_HWDATA_0_iv_17_920_0_0, 
        un1_hready_2, N_4827, N_450, N_228, d_HWRITE_0_sqmuxa_4, 
        un1_state_30, N_582, N_4874, N_683_2, N_4873, N_4556_1, 
        N_682_2, N_686_2, N_96, N_182_1, \un1_state_39\, 
        \un1_state_46_0\, \state_m2_e_1\, 
        d_HWDATA_0_iv_6_1388_5_0, d_HWDATA_0_iv_2_1532_5_0, 
        d_HWDATA_0_iv_1_1568_0_1, N_929, N_444, N_4764, N_4837, 
        N_453, N_285, N_286, N_287, N_296, \ins2_i_m[17]\, N_4387, 
        \ins2_m[23]\, \ins2_m[19]\, \ins2_m[26]\, \ins2_m[25]\, 
        \ins2_m[28]\, \ins2_m[20]\, \ins2_m[2]\, N_4445, N_4514, 
        N_4524, N_4759, \ins2_m[9]\, N_4854, N_4857, N_4519, 
        N_411_2, N_212, \d_count_0_0_0[1]\, 
        \d_HADDR_0_iv_0_0[0]_net_1\, \d_HADDR_0_iv_0[2]_net_1\, 
        \d_HADDR_0_iv_0_0[17]_net_1\, \d_HADDR_0_iv_0[9]_net_1\, 
        \d_HADDR_0_iv_0_0[5]_net_1\, \d_HADDR_0_iv_0[28]_net_1\, 
        \d_HADDR_0_iv_0[23]_net_1\, \d_HADDR_0_iv_0[25]_net_1\, 
        \d_HADDR_0_iv_0[19]_net_1\, \d_HADDR_0_iv_0[26]_net_1\, 
        \d_HADDR_0_iv_0_0[18]_net_1\, 
        \d_HADDR_0_iv_0_0[16]_net_1\, 
        \d_HADDR_0_iv_0_0[21]_net_1\, \d_HADDR_0_iv_0[20]_net_1\, 
        \d_HADDR_0_iv_0_0[12]_net_1\, 
        \d_HADDR_0_iv_0_0[10]_net_1\, \state_m3_i_7\, 
        \un1_state_46_1\, \d_count_i_2[0]\, \un1_state_44_0_12\, 
        \un1_d_HWRITE_0_sqmuxa_5_i_0_2\, 
        \un1_d_HWRITE_0_sqmuxa_5_i_0_0\, \un1_state_42_0_0_3\, 
        \d_count_0_a2_1_c_1[1]\, \state_m2_e_2\, 
        \d_count_0_o3_3_1[1]\, N_186, 
        \state_ns_i_0_a2_3_d_0[1]_net_1\, \d_HWDATA_0_sqmuxa_2\, 
        N_4856, \state_m3_i_8\, N_148, \un1_state_46_3\, 
        \d_count_0_2[1]\, \state_m3_i_a3\, 
        \d_HADDR_0_iv_2[2]_net_1\, \d_HADDR_0_iv_0_2[17]_net_1\, 
        \d_HADDR_0_iv_2[9]_net_1\, \d_HADDR_0_iv_0_2[5]_net_1\, 
        \d_HADDR_0_iv_2[28]_net_1\, \d_HADDR_0_iv_2[23]_net_1\, 
        \d_HADDR_0_iv_2[25]_net_1\, \d_HADDR_0_iv_2[19]_net_1\, 
        \d_HADDR_0_iv_2[26]_net_1\, \d_HADDR_0_iv_0_2[18]_net_1\, 
        \d_HADDR_0_iv_0_2[16]_net_1\, 
        \d_HADDR_0_iv_0_2[21]_net_1\, \d_HADDR_0_iv_2[20]_net_1\, 
        \d_HADDR_0_iv_0_2[12]_net_1\, 
        \d_HADDR_0_iv_0_2[10]_net_1\ : std_logic;

begin 

    ConfigMaster_0_M_HADDR(31) <= \ConfigMaster_0_M_HADDR[31]\;
    ConfigMaster_0_M_HADDR(30) <= \ConfigMaster_0_M_HADDR[30]\;
    ConfigMaster_0_M_HADDR(29) <= \ConfigMaster_0_M_HADDR[29]\;
    ConfigMaster_0_M_HADDR(28) <= \ConfigMaster_0_M_HADDR[28]\;
    ConfigMaster_0_M_HADDR(27) <= \ConfigMaster_0_M_HADDR[27]\;
    ConfigMaster_0_M_HADDR(26) <= \ConfigMaster_0_M_HADDR[26]\;
    ConfigMaster_0_M_HADDR(25) <= \ConfigMaster_0_M_HADDR[25]\;
    ConfigMaster_0_M_HADDR(24) <= \ConfigMaster_0_M_HADDR[24]\;
    ConfigMaster_0_M_HADDR(23) <= \ConfigMaster_0_M_HADDR[23]\;
    ConfigMaster_0_M_HADDR(22) <= \ConfigMaster_0_M_HADDR[22]\;
    ConfigMaster_0_M_HADDR(21) <= \ConfigMaster_0_M_HADDR[21]\;
    ConfigMaster_0_M_HADDR(20) <= \ConfigMaster_0_M_HADDR[20]\;
    ConfigMaster_0_M_HADDR(19) <= \ConfigMaster_0_M_HADDR[19]\;
    ConfigMaster_0_M_HADDR(18) <= \ConfigMaster_0_M_HADDR[18]\;
    ConfigMaster_0_M_HADDR(17) <= \ConfigMaster_0_M_HADDR[17]\;
    ConfigMaster_0_M_HADDR(16) <= \ConfigMaster_0_M_HADDR[16]\;
    ConfigMaster_0_M_HADDR(15) <= \ConfigMaster_0_M_HADDR[15]\;
    ConfigMaster_0_M_HADDR(14) <= \ConfigMaster_0_M_HADDR[14]\;
    ConfigMaster_0_M_HADDR(13) <= \ConfigMaster_0_M_HADDR[13]\;
    ConfigMaster_0_M_HADDR(12) <= \ConfigMaster_0_M_HADDR[12]\;
    ConfigMaster_0_M_HADDR(11) <= \ConfigMaster_0_M_HADDR[11]\;
    ConfigMaster_0_M_HADDR(10) <= \ConfigMaster_0_M_HADDR[10]\;
    ConfigMaster_0_M_HADDR(9) <= \ConfigMaster_0_M_HADDR[9]\;
    ConfigMaster_0_M_HADDR(8) <= \ConfigMaster_0_M_HADDR[8]\;
    ConfigMaster_0_M_HADDR(7) <= \ConfigMaster_0_M_HADDR[7]\;
    ConfigMaster_0_M_HADDR(6) <= \ConfigMaster_0_M_HADDR[6]\;
    ConfigMaster_0_M_HADDR(5) <= \ConfigMaster_0_M_HADDR[5]\;
    ConfigMaster_0_M_HADDR(4) <= \ConfigMaster_0_M_HADDR[4]\;
    ConfigMaster_0_M_HADDR(3) <= \ConfigMaster_0_M_HADDR[3]\;
    ConfigMaster_0_M_HADDR(2) <= \ConfigMaster_0_M_HADDR[2]\;
    ConfigMaster_0_M_HADDR(1) <= \ConfigMaster_0_M_HADDR[1]\;
    ConfigMaster_0_M_HADDR(0) <= \ConfigMaster_0_M_HADDR[0]\;

    \d_HADDR_0_iv_0[2]\ : CFG4
      generic map(INIT => x"5D0C")

      port map(A => \ConfigMaster_0_M_HADDR[2]\, B => 
        \haddr_write[2]_net_1\, C => N_4874, D => un1_state_30, Y
         => \d_HADDR_0_iv_0[2]_net_1\);
    
    un1_rdata_0_I_50_i_0_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[22]_net_1\, B => \rdata[22]_net_1\, 
        C => \mask[22]_net_1\, Y => N_359_i);
    
    un1_d_HWRITE_0_sqmuxa_5_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \state[11]_net_1\, B => \state[10]_net_1\, C
         => N_259, Y => N_137);
    
    un7_hready_2_RNI3VJ11 : CFG2
      generic map(INIT => x"8")

      port map(A => N_591, B => N_251, Y => N_512_1);
    
    un1_rdata_0_I_98_i_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[25]_net_1\, B => \rdata[25]_net_1\, 
        C => \mask[25]_net_1\, Y => N_327_i);
    
    \HWDATA_int[15]\ : SLE
      port map(D => \HWDATA_int_RNO[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(15));
    
    un1_state_39_3 : CFG2
      generic map(INIT => x"E")

      port map(A => \state[13]_net_1\, B => \state[18]_net_1\, Y
         => \un1_state_39_3\);
    
    \HWDATA_int_RNO_0[13]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[13]_net_1\, D => \rdata[29]_net_1\, Y => 
        d_HWDATA_0_iv_17_920_0_0);
    
    \d_HADDR_0_iv_0[14]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => un13_d_haddr_1_s_12_S, B => \state_ns[0]\, C
         => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0[14]_net_1\);
    
    \ins2[5]\ : SLE
      port map(D => \d_ins2[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[5]_net_1\);
    
    \HWDATA_int_RNO_2[26]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[22]_net_1\, B => \rdata[10]_net_1\, C
         => N_276, D => \count[1]_net_1\, Y => N_4577);
    
    \haddr_fetch[9]\ : SLE
      port map(D => N_4418_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[9]_net_1\);
    
    \HWDATA_int_RNO_0[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_270, C => 
        \acc[1]_net_1\, D => \rdata[1]_net_1\, Y => 
        d_HWDATA_0_iv_29_425_0_0);
    
    \state[23]\ : SLE
      port map(D => \state_ns[5]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[23]_net_1\);
    
    \haddr_fetch[22]\ : SLE
      port map(D => N_4722_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[22]_net_1\);
    
    un1_rdata_0_I_28 : CFG3
      generic map(INIT => x"6A")

      port map(A => \expected[7]_net_1\, B => \rdata[7]_net_1\, C
         => \mask[7]_net_1\, Y => un1_rdata_0_N_57);
    
    \d_HADDR_0_iv_0_0[5]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_3_S, B => 
        \haddr_write[5]_net_1\, C => N_4874, D => un1_state_30, Y
         => \d_HADDR_0_iv_0_0[5]_net_1\);
    
    un1_state_42_0_0 : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \ins1[31]_net_1\, B => N_182_1, C => 
        \un1_state_42_0_0_3\, D => N_929, Y => \un1_state_42_0_0\);
    
    \HADDR_int[15]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[15]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[15]\);
    
    \HWDATA_int_RNO_0[4]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_270, C => 
        \acc[4]_net_1\, D => \rdata[4]_net_1\, Y => 
        d_HWDATA_0_iv_26_560_0_0);
    
    \haddr_write[7]\ : SLE
      port map(D => un46_d_haddr_cry_7_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[7]_net_1\);
    
    un1_state_44_0_o2_0 : CFG4
      generic map(INIT => x"FFFD")

      port map(A => N_837, B => \state[23]_net_1\, C => N_4814, D
         => N_117, Y => N_4827);
    
    d_HWRITE_0_sqmuxa_2_0_a3 : CFG3
      generic map(INIT => x"40")

      port map(A => N_290, B => d_N_3_mux_0, C => 
        \d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0\, Y => 
        d_HWRITE_0_sqmuxa_2);
    
    \state_ns_i_a2_10_i_o2[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \state[10]_net_1\, B => \state[11]_net_1\, Y
         => N_138);
    
    \HWDATA_int[9]\ : SLE
      port map(D => \HWDATA_int_RNO[9]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(9));
    
    \un7_iv_0_a1_0[14]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_252, B => \state_21_rep1\, Y => 
        \un7_iv_0_a1_0[14]_net_1\);
    
    \HADDR_int_fast[0]\ : SLE
      port map(D => \d_HADDR_fast[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \HADDR_int_fast[0]_net_1\);
    
    \expected[4]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(4), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[4]_net_1\);
    
    \state[25]\ : SLE
      port map(D => N_70_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[25]_net_1\);
    
    \state[28]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[28]_net_1\);
    
    \d_HADDR_0_iv_1_0[29]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_1[29]_net_1\, B => 
        \haddr_fetch[29]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1_0[29]_net_1\);
    
    \ins1_RNINCALRA[14]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[14]_net_1\, B => N_78, C => N_164, 
        D => \ins1[14]_net_1\, FCI => d_bytecount_i_m2_cry_13, S
         => N_116, Y => OPEN, FCO => d_bytecount_i_m2_cry_14);
    
    \expected[5]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(5), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[5]_net_1\);
    
    \haddr_fetch[4]\ : SLE
      port map(D => N_2921_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[4]_net_1\);
    
    un46_d_haddr_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[10]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_9\, S => un46_d_haddr_cry_10_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_10\);
    
    \d_HADDR_0_iv_0[18]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[18]_net_1\, C => 
        \haddr_fetch[18]_net_1\, Y => \d_HADDR[18]\);
    
    \ins1_RNIE4ISO[0]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[0]_net_1\, B => N_78, C => N_166, 
        D => \ins1[0]_net_1\, FCI => GND_net_1, S => OPEN, Y => 
        \ins1_RNIE4ISO_Y[0]\, FCO => d_bytecount_i_m2_cry_0);
    
    \HWDATA_int_RNO_0[22]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \state[10]_net_1\, B => N_4653, C => 
        \acc[22]_net_1\, Y => d_HWDATA_0_iv_8_1298_1_0);
    
    \d_acc[12]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1149, C => 
        \ins2[12]_net_1\, D => \acc[12]_net_1\, Y => 
        \d_acc[12]_net_1\);
    
    \rdata_RNI95Q62[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \rdata[26]_net_1\, B => \rdata[10]_net_1\, C
         => N_655, D => N_600, Y => N_286);
    
    \ins1_RNIVQ38Q7[10]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[10]_net_1\, B => N_78, C => N_164, 
        D => \ins1[10]_net_1\, FCI => d_bytecount_i_m2_cry_9, S
         => N_4339, Y => OPEN, FCO => d_bytecount_i_m2_cry_10);
    
    \d_HADDR_0_iv_2[11]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[11]_net_1\, B => 
        \ins2[11]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_2[11]_net_1\);
    
    un1_state_42_0_o2_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[24]_net_1\, B => \state[23]_net_1\, C
         => \state[14]_net_1\, D => \state[11]_net_1\, Y => N_136);
    
    \haddr_write[24]\ : SLE
      port map(D => un46_d_haddr_cry_24_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[24]_net_1\);
    
    un1_state_31_i_i_a2_0_d_0_0_1 : CFG4
      generic map(INIT => x"0001")

      port map(A => N_98, B => N_25, C => 
        defSlaveSMNextState_m_0_3_1, D => 
        defSlaveSMNextState_m_0_2, Y => 
        \un1_state_31_i_i_a2_0_d_0_0_1\);
    
    \mask[16]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(16), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[16]_net_1\);
    
    un1_state_44_0_a3_3 : CFG4
      generic map(INIT => x"E400")

      port map(A => N_109_i, B => un1_hready_2, C => 
        \ins1[31]_net_1\, D => \state[21]_net_1\, Y => N_4856);
    
    \ins1_RNIACDJI8[11]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[11]_net_1\, B => N_78, C => N_164, 
        D => \ins1[11]_net_1\, FCI => d_bytecount_i_m2_cry_10, S
         => N_4340, Y => OPEN, FCO => d_bytecount_i_m2_cry_11);
    
    \d_HADDR_0_iv_0_2[10]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_10_S, B => 
        \d_HADDR_0_iv_0_0[10]_net_1\, C => N_4519, D => N_247, Y
         => \d_HADDR_0_iv_0_2[10]_net_1\);
    
    \HWDATA_int_RNO_1[26]\ : CFG4
      generic map(INIT => x"B3A0")

      port map(A => \state[10]_net_1\, B => N_263, C => 
        \acc[26]_net_1\, D => \rdata[10]_net_1\, Y => 
        d_HWDATA_0_iv_4_1460_5_0);
    
    \HADDR_int[9]\ : SLE
      port map(D => \d_HADDR[9]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[9]\);
    
    \expected[25]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(25), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[25]_net_1\);
    
    \ins1_RNI6L0A3A[13]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[13]_net_1\, B => N_78, C => N_164, 
        D => \ins1[13]_net_1\, FCI => d_bytecount_i_m2_cry_12, S
         => N_4341, Y => OPEN, FCO => d_bytecount_i_m2_cry_13);
    
    \d_HADDR_0_iv[26]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[26]_net_1\, C => \haddr_fetch[26]_net_1\, 
        Y => \d_HADDR[26]\);
    
    \ins1_RNIUC04_1[22]\ : CFG4
      generic map(INIT => x"0110")

      port map(A => \ins1[23]_net_1\, B => \ins1[22]_net_1\, C
         => \ins1[21]_net_1\, D => \ins1[20]_net_1\, Y => N_290);
    
    un46_d_haddr_cry_24 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[24]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_23\, S => un46_d_haddr_cry_24_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_24\);
    
    \d_acc_0[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[2]_net_1\, B => \ins2[2]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(2), D => \state[8]_net_1\, Y => 
        N_1139);
    
    \state_ns_0_fast[7]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \state_fast[21]_net_1\, B => 
        d_state_1_sqmuxa_1_i_0, C => N_109_i, D => N_101, Y => 
        \state_ns_fast[7]\);
    
    \acc[27]\ : SLE
      port map(D => \d_acc[27]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[27]_net_1\);
    
    \ins2[20]\ : SLE
      port map(D => \d_ins2[20]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[20]_net_1\);
    
    \rdata_RNIR09F[15]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \state[21]_net_1\, B => \count[1]_net_1\, C
         => \rdata[15]_net_1\, Y => N_2066);
    
    \ins1[5]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(5), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[5]_net_1\);
    
    \d_acc_0[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[1]_net_1\, B => \ins2[1]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(1), D => \state[8]_net_1\, Y => 
        N_1138);
    
    \ins1_RNIT0FT86[8]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[8]_net_1\, B => N_78, C => N_164, 
        D => \ins1[8]_net_1\, FCI => d_bytecount_i_m2_cry_7, S
         => N_4337, Y => OPEN, FCO => d_bytecount_i_m2_cry_8);
    
    \rdata_RNI68SG[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \rdata[0]_net_1\, B => \count[1]_net_1\, C
         => N_249, Y => N_465);
    
    un1_state_44_0_a3_1 : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \state[25]_net_1\, B => \ins1[25]_net_1\, C
         => N_198, D => HREADY_i_3, Y => N_4854);
    
    \ins1[29]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(29), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[29]_net_1\);
    
    \rdata_RNINB9J[13]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => \rdata[13]_net_1\, B => N_263, C => N_249, Y
         => N_4885);
    
    \d_HADDR_0_iv_0_0[12]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_10_S, B => 
        \haddr_write[12]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[12]_net_1\);
    
    \ins2[8]\ : SLE
      port map(D => \d_ins2[8]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[8]_net_1\);
    
    \d_acc_0[14]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[14]_net_1\, B => \ins2[14]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(14), D => \state[8]_net_1\, Y => 
        N_1151);
    
    \expected[18]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(18), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[18]_net_1\);
    
    \haddr_write[21]\ : SLE
      port map(D => un46_d_haddr_cry_21_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[21]_net_1\);
    
    \state[17]\ : SLE
      port map(D => \state_ns[11]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[17]_net_1\);
    
    \d_ins2[26]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(26), B => un28_opcode, 
        Y => \d_ins2[26]_net_1\);
    
    \state[6]\ : SLE
      port map(D => \state_ns[22]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[6]_net_1\);
    
    \d_HADDR_0_iv_0_0_1[24]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => N_481, B => \haddr_fetch[24]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_0_0_1[24]_net_1\);
    
    \HWDATA_int[23]\ : SLE
      port map(D => \HWDATA_int_RNO[23]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(23));
    
    \HADDR_int[7]\ : SLE
      port map(D => \d_HADDR[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[7]\);
    
    \d_HADDR_0_iv_0[25]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_23_S, B => 
        \haddr_write[25]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[25]_net_1\);
    
    \expected[21]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(21), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[21]_net_1\);
    
    \acc[1]\ : SLE
      port map(D => \d_acc[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[1]_net_1\);
    
    \haddr_write[31]\ : SLE
      port map(D => un46_d_haddr_s_31_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[31]_net_1\);
    
    \d_ins2[23]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(23), B => un28_opcode, 
        Y => \d_ins2[23]_net_1\);
    
    \count_RNIGI2A_0[1]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \count[1]_net_1\, B => \state[21]_net_1\, Y
         => N_272);
    
    \state_RNIBKIN[22]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \state[22]_net_1\, B => \count[0]_net_1\, C
         => \state[21]_net_1\, D => N_249, Y => N_262);
    
    \HWDATA_int_RNO_0[31]\ : CFG4
      generic map(INIT => x"3133")

      port map(A => N_276, B => d_HWDATA_0_iv_1640_2, C => 
        \count[1]_net_1\, D => N_2573_1, Y => 
        d_HWDATA_0_iv_1640_1);
    
    un1_hready_2_0_a2_RNI1ABB : CFG2
      generic map(INIT => x"D")

      port map(A => N_252, B => N_4912, Y => 
        d_state_1_sqmuxa_1_i_0);
    
    \state_ns_0_a3_2_0[8]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \state[4]_net_1\, B => N_133, C => 
        \state[3]_net_1\, D => \ins1[31]_net_1\, Y => 
        \state_ns_0_a3_2[8]_net_1\);
    
    \d_HADDR_0_iv_RNO[22]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => un13_d_haddr_1_cry_20_S, B => 
        \un1_state_30_0_0\, C => N_4814, Y => 
        \un13_d_haddr_1_m[22]\);
    
    un1_rdata_0_I_45 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[23]_net_1\, B => N_359_i, C => 
        \expected[23]_net_1\, D => \mask[23]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[10]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[11]\);
    
    \mask[17]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(17), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[17]_net_1\);
    
    un1_rdata_0_I_33 : ARI1
      generic map(INIT => x"40095")

      port map(A => un1_rdata_0_N_53, B => \expected[21]_net_1\, 
        C => \mask[21]_net_1\, D => \rdata[21]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[9]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[10]\);
    
    \acc[14]\ : SLE
      port map(D => \d_acc[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[14]_net_1\);
    
    un1_state_39_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \un1_state_39_1_0_a3_0_1\, B => 
        \un1_state_39_3\, C => N_200, D => N_80, Y => 
        \un1_state_39_1\);
    
    \expected[31]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(31), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[31]_net_1\);
    
    un1_rdata_0_I_68_i_0_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[10]_net_1\, B => \rdata[10]_net_1\, 
        C => \mask[10]_net_1\, Y => N_351_i);
    
    un13_d_haddr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[3]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un13_d_haddr_1_s_1_172_FCO, S => un13_d_haddr_1_cry_1_S, 
        Y => OPEN, FCO => \un13_d_haddr_1_cry_1\);
    
    \haddr_fetch[17]\ : SLE
      port map(D => N_4403_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[17]_net_1\);
    
    \bytecount[12]\ : SLE
      port map(D => N_50_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[12]_net_1\);
    
    \state_fast_RNIDMVC[21]\ : CFG4
      generic map(INIT => x"111D")

      port map(A => \state[22]_net_1\, B => 
        \state_fast[21]_net_1\, C => \count[1]_net_1\, D => 
        \count[0]_net_1\, Y => un1_state_31_i_i_o2_0);
    
    \ins1_RNIMBQS17[9]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[9]_net_1\, B => N_78, C => N_164, 
        D => \ins1[9]_net_1\, FCI => d_bytecount_i_m2_cry_8, S
         => N_4338, Y => OPEN, FCO => d_bytecount_i_m2_cry_9);
    
    \HSIZE_int[0]\ : SLE
      port map(D => N_415, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_34_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HSIZE(0));
    
    \d_HADDR_0_iv_0_1[13]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_0_0[13]_net_1\, B => 
        \haddr_fetch[13]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_0_1[13]_net_1\);
    
    \bytecount[1]\ : SLE
      port map(D => \d_bytecount[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[1]_net_1\);
    
    un46_d_haddr_cry_25 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[25]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_24\, S => un46_d_haddr_cry_25_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_25\);
    
    \expected[9]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(9), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[9]_net_1\);
    
    \d_acc_1[3]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[3]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(3), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[3]\);
    
    \envm_busy[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_14_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \envm_busy[1]_net_1\);
    
    \HWDATA_int_RNO_1[15]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \rdata[31]_net_1\, B => \state[21]_net_1\, C
         => N_4879, D => d_HWDATA_0_iv_15_992_2, Y => 
        d_HWDATA_0_iv_15_992_4);
    
    \HWDATA_int_RNO_0[23]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_601, C => 
        \acc[23]_net_1\, D => \rdata[7]_net_1\, Y => 
        d_HWDATA_0_iv_7_1343_1_0);
    
    \acc[9]\ : SLE
      port map(D => \d_acc[9]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[9]_net_1\);
    
    \HADDR_int_RNO_1[15]\ : CFG4
      generic map(INIT => x"4445")

      port map(A => \d_HADDR_0_iv_1[15]_net_1\, B => 
        \haddr_fetch[15]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => \d_HADDR_0_iv_i_1[15]\);
    
    \HWDATA_int[18]\ : SLE
      port map(D => \HWDATA_int_RNO[18]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(18));
    
    \HWDATA_int[2]\ : SLE
      port map(D => \HWDATA_int_RNO[2]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(2));
    
    \bytecount[5]\ : SLE
      port map(D => N_36_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[5]_net_1\);
    
    un1_state_42_0_o2 : CFG2
      generic map(INIT => x"7")

      port map(A => d_state61_li, B => \ins1[31]_net_1\, Y => 
        N_125);
    
    \haddr_fetch_RNO[17]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_15_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[17]\, D => N_4812, Y => 
        N_4403_i_0);
    
    un46_d_haddr_cry_29 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[29]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_28\, S => un46_d_haddr_cry_29_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_29\);
    
    \d_HADDR_0_iv_0_2[3]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => \haddr_write[3]_net_1\, B => \ins2[3]_net_1\, 
        C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_0_2[3]_net_1\);
    
    \d_HADDR_0_iv_2[26]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_26_S, B => 
        \d_HADDR_0_iv_0[26]_net_1\, C => \ins2_m[26]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[26]_net_1\);
    
    \rdata[19]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(19), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[19]_net_1\);
    
    \HWDATA_int[8]\ : SLE
      port map(D => \HWDATA_int_RNO[8]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(8));
    
    \d_HADDR_0_iv_2[28]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_28_S, B => 
        \d_HADDR_0_iv_0[28]_net_1\, C => \ins2_m[28]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[28]_net_1\);
    
    un46_d_haddr_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[11]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_10\, S => un46_d_haddr_cry_11_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_11\);
    
    \HWDATA_int_RNO_3[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \state[10]_net_1\, B => N_2066, C => 
        \acc[15]_net_1\, Y => d_HWDATA_0_iv_15_992_0);
    
    un13_d_haddr_1_cry_19 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[21]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_18\, S => un13_d_haddr_1_cry_19_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_19\);
    
    \HWDATA_int_RNO[12]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_18_884_6_0, B => N_686_2, C => 
        \rdata[12]_net_1\, D => N_264, Y => 
        \HWDATA_int_RNO[12]_net_1\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o3_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_109_i, B => un1_state_31_i_i_a2_0_d_1_0_1, 
        C => N_4912, D => un1_d_HWRITE_1_sqmuxa_2_i_o3_1_0, Y => 
        un1_d_HWRITE_1_sqmuxa_2_i_o3_1_2);
    
    d_haddr_fetch_2_sqmuxa_0 : CFG2
      generic map(INIT => x"4")

      port map(A => N_198, B => \state[25]_net_1\, Y => 
        \d_haddr_fetch_2_sqmuxa_0\);
    
    \d_HADDR_0_iv_0[20]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_18_S, B => 
        \haddr_write[20]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[20]_net_1\);
    
    un13_d_haddr_1_cry_27_5 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[14]\, B => 
        \ConfigMaster_0_M_HADDR[11]\, C => 
        \ConfigMaster_0_M_HADDR[12]\, D => 
        \ConfigMaster_0_M_HADDR[13]\, FCI => 
        un13_d_haddr_1_cry_27_3_FCO, S => OPEN, Y => OPEN, FCO
         => un13_d_haddr_1_cry_27_5_FCO);
    
    \rdata_RNI02TD2[25]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => N_585, B => \rdata[25]_net_1\, C => N_582, D
         => N_257, Y => N_296);
    
    \ins2[19]\ : SLE
      port map(D => \d_ins2[19]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[19]_net_1\);
    
    \ins2[26]\ : SLE
      port map(D => \d_ins2[26]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[26]_net_1\);
    
    \d_bytecount[1]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_1102, B => \state[21]_net_1\, C => N_109_i, 
        Y => \d_bytecount[1]_net_1\);
    
    \state[2]\ : SLE
      port map(D => N_14_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[2]_net_1\);
    
    un1_rdata_0_I_9 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[29]_net_1\, B => N_355_i, C => 
        \expected[29]_net_1\, D => \mask[29]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[13]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[14]\);
    
    \rdata_RNIB7Q62[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \rdata[27]_net_1\, B => \rdata[11]_net_1\, C
         => N_655, D => N_600, Y => N_288);
    
    \count_RNINH9E1[0]\ : CFG4
      generic map(INIT => x"FBF3")

      port map(A => N_272, B => \count[0]_net_1\, C => 
        d_HWDATA_0_iv_14_1028_0_a2_i_1, D => N_317, Y => N_178);
    
    \haddr_write[26]\ : SLE
      port map(D => un46_d_haddr_cry_26_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[26]_net_1\);
    
    \rdata[27]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(27), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[27]_net_1\);
    
    \d_HADDR_0_iv_1_0[27]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_1[27]_net_1\, B => 
        \haddr_fetch[27]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1_0[27]_net_1\);
    
    \HWDATA_int_RNO[22]\ : CFG4
      generic map(INIT => x"FBBB")

      port map(A => d_HWDATA_0_iv_8_1298_1_0, B => N_4891, C => 
        \rdata[22]_net_1\, D => N_4625, Y => 
        \HWDATA_int_RNO[22]_net_1\);
    
    un46_d_haddr_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[6]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_5\, S => un46_d_haddr_cry_6_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_6\);
    
    un1_d_HWRITE_0_sqmuxa_1_0_a3_i_1 : CFG4
      generic map(INIT => x"DFCF")

      port map(A => N_266, B => N_272, C => N_276, D => 
        d_N_3_mux_0, Y => \un1_d_HWRITE_0_sqmuxa_1_0_a3_i_1\);
    
    \d_HADDR_0_iv_0[19]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_17_S, B => 
        \haddr_write[19]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[19]_net_1\);
    
    \HADDR_int[8]\ : SLE
      port map(D => \d_HADDR[8]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[8]\);
    
    \ins1[20]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(20), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[20]_net_1\);
    
    \state[19]\ : SLE
      port map(D => \state_ns[9]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[19]_net_1\);
    
    d_HTRANS_0_sqmuxa_4_1_1_o3_1_RNIK29J2 : CFG4
      generic map(INIT => x"0800")

      port map(A => \un12_size_2_0_4\, B => d_m1_e_1_1, C => 
        \d_HTRANS_0_sqmuxa_4_1_1_o3_1\, D => \un12_size_2_0_5\, Y
         => d_N_3_mux_0);
    
    \d_HADDR_0_iv_0_a2_3[10]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[10]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4519);
    
    \HWDATA_int[19]\ : SLE
      port map(D => \HWDATA_int_RNO[19]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(19));
    
    un1_hready_2_0_a2_RNIQ8TL : CFG4
      generic map(INIT => x"B1BB")

      port map(A => \state_21_rep1\, B => \state[22]_net_1\, C
         => N_4912, D => N_252, Y => 
        un1_state_31_i_i_a2_0_d_0_0_0);
    
    \mask[25]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(25), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[25]_net_1\);
    
    \ins2[31]\ : SLE
      port map(D => \d_ins2[31]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[31]_net_1\);
    
    un13_d_haddr_1_cry_27_3 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[10]\, B => 
        \ConfigMaster_0_M_HADDR[7]\, C => 
        \ConfigMaster_0_M_HADDR[8]\, D => 
        \ConfigMaster_0_M_HADDR[9]\, FCI => 
        un13_d_haddr_1_cry_27_1_FCO, S => OPEN, Y => OPEN, FCO
         => un13_d_haddr_1_cry_27_3_FCO);
    
    state_21_rep1_RNIEVN4O : CFG4
      generic map(INIT => x"FEEE")

      port map(A => un1_state_31_i_i_a2_0_d_1_sx_0, B => 
        un1_state_31_i_i_a2_0_d_1_0_sx, C => \state_21_rep1\, D
         => defSlaveSMNextState_m_0_3, Y => N_166);
    
    \d_HADDR_0_iv[4]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_2[4]_net_1\, B => 
        un46_d_haddr_cry_4_S, C => \d_HADDR_0_iv_1[4]_net_1\, D
         => N_247, Y => \d_HADDR[4]\);
    
    \d_bytecount[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_1104, B => \state[21]_net_1\, C => N_109_i, 
        Y => \d_bytecount[3]_net_1\);
    
    \d_acc_0[15]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[15]_net_1\, B => \ins2[15]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(15), D => \state[8]_net_1\, Y => 
        N_1152);
    
    \d_acc[26]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1163, C => 
        \ins2[26]_net_1\, D => \acc[26]_net_1\, Y => 
        \d_acc[26]_net_1\);
    
    \HWDATA_int_RNO_1[31]\ : CFG4
      generic map(INIT => x"DDFD")

      port map(A => d_HWDATA_0_iv_1640_2_1, B => N_2579, C => 
        d_HWDATA_0_iv_1640_a8_3_0, D => N_252, Y => 
        d_HWDATA_0_iv_1640_2);
    
    \haddr_fetch[31]\ : SLE
      port map(D => N_4366_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[31]_net_1\);
    
    \rdata_RNID0SC[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \count[1]_net_1\, B => \rdata[5]_net_1\, Y
         => N_4539);
    
    \rdata_RNINCAJ[23]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[21]_net_1\, B => N_249, C => 
        \rdata[23]_net_1\, D => \count[0]_net_1\, Y => N_2579);
    
    \bytecount_RNO[2]\ : CFG3
      generic map(INIT => x"70")

      port map(A => \state[21]_net_1\, B => N_109_i, C => N_104, 
        Y => N_32_i_0);
    
    un1_rdata_0_I_75 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[17]_net_1\, B => N_323_i, C => 
        \expected[17]_net_1\, D => \mask[17]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[7]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[8]\);
    
    un13_d_haddr_1_cry_26 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[28]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_25\, S => un13_d_haddr_1_cry_26_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_26\);
    
    \expected[28]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(28), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[28]_net_1\);
    
    \acc[30]\ : SLE
      port map(D => \d_acc[30]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[30]_net_1\);
    
    un1_rdata_0_I_63 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[11]_net_1\, B => N_351_i, C => 
        \expected[11]_net_1\, D => \mask[11]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[4]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[5]\);
    
    \acc[2]\ : SLE
      port map(D => \d_acc[2]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[2]_net_1\);
    
    \HWDATA_int_RNO_4[15]\ : CFG4
      generic map(INIT => x"4500")

      port map(A => \count[1]_net_1\, B => \count[0]_net_1\, C
         => N_249, D => N_2573_1, Y => N_2063);
    
    \haddr_write[18]\ : SLE
      port map(D => un46_d_haddr_cry_18_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[18]_net_1\);
    
    \haddr_fetch[30]\ : SLE
      port map(D => N_17_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[30]_net_1\);
    
    \HWDATA_int_RNO_2[25]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[22]_net_1\, B => \rdata[9]_net_1\, C
         => N_276, D => \count[1]_net_1\, Y => N_2399);
    
    \HADDR_int[21]\ : SLE
      port map(D => \d_HADDR[21]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[21]\);
    
    un1_state_34_0_0 : CFG3
      generic map(INIT => x"AE")

      port map(A => N_929, B => \state[24]_net_1\, C => 
        HREADY_i_3, Y => \un1_state_34_0_0\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bytecount_RNO[9]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4338, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_44_i_0);
    
    \acc[23]\ : SLE
      port map(D => \d_acc[23]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[23]_net_1\);
    
    \d_acc_0[12]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[12]_net_1\, B => \ins2[12]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(12), D => \state[8]_net_1\, Y => 
        N_1149);
    
    \d_HADDR_0_iv_2[6]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => \haddr_write[6]_net_1\, B => \ins2[6]_net_1\, 
        C => N_4873, D => N_4874, Y => \d_HADDR_0_iv_2[6]_net_1\);
    
    \HWDATA_int_RNO[15]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_2060, B => N_2579, C => 
        d_HWDATA_0_iv_15_992_4, D => N_2061, Y => 
        \HWDATA_int_RNO[15]_net_1\);
    
    d_HWRITE_0_sqmuxa_4_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => \d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0\, B => 
        \state[22]_net_1\, C => d_N_3_mux_0, D => N_249, Y => 
        N_402);
    
    \un7_iv_1[14]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => defSlaveSMNextState_i_a2_0_RNI3J724_2, B => 
        N_252, C => defSlaveSMNextState_m_0_3, D => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, Y => 
        \un7_iv_1[14]_net_1\);
    
    \state[16]\ : SLE
      port map(D => N_480, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[16]_net_1\);
    
    un1_state_44_0_a3_4 : CFG3
      generic map(INIT => x"08")

      port map(A => \ins1[31]_net_1\, B => N_117, C => HREADY_i_3, 
        Y => N_4857);
    
    \d_HADDR_0_iv_0_a2_3[12]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[12]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4445);
    
    \mask[9]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(9), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[9]_net_1\);
    
    \rdata_RNI8AMI[21]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_4539, B => N_4541, Y => N_4472);
    
    \d_HADDR_0_iv_0_0[30]\ : CFG4
      generic map(INIT => x"DDDC")

      port map(A => un13_d_haddr_1_cry_28_S, B => \state_ns[0]\, 
        C => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0_0[30]_net_1\);
    
    \HWDATA_int_RNO[25]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => d_HWDATA_0_iv_5_1424_1, B => N_2380_3, C => 
        N_2400, D => N_2399, Y => \HWDATA_int_RNO[25]_net_1\);
    
    \HWDATA_int_RNO[2]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_28_470_3_0, B => N_286, C => 
        \rdata[18]_net_1\, D => N_271, Y => 
        \HWDATA_int_RNO[2]_net_1\);
    
    \d_acc_1_0_0[24]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[24]_net_1\, B => \acc[24]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0_0[24]_net_1\);
    
    \pause_count_RNO[4]\ : CFG4
      generic map(INIT => x"00CE")

      port map(A => \pause_count[3]_net_1\, B => 
        \pause_count[4]_net_1\, C => N_4811, D => N_3400, Y => 
        N_4809_i_0);
    
    \ins2[10]\ : SLE
      port map(D => \d_ins2[10]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[10]_net_1\);
    
    \HWDATA_int_RNO_0[9]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[9]_net_1\, D => \rdata[25]_net_1\, Y => 
        d_HWDATA_0_iv_21_776_6_0);
    
    \d_acc_1_0[5]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[5]_net_1\, B => \acc[5]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[5]_net_1\);
    
    \haddr_write[29]\ : SLE
      port map(D => un46_d_haddr_cry_29_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[29]_net_1\);
    
    \state_ns_i_a2_13_0_a3_8[1]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_117, B => 
        \state_ns_i_a2_13_0_a3_5[1]_net_1\, C => N_136, D => 
        N_200, Y => \state_ns_i_a2_13_0_a3_8[1]_net_1\);
    
    \haddr_fetch_RNO[12]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_10_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[12]\, D => N_4812, Y => 
        N_4402_i_0);
    
    un1_state_44_0_9 : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \busy\, B => \state[1]_net_1\, C => 
        \un1_state_44_0_4\, D => \un1_state_44_0_8\, Y => 
        \un1_state_44_0_9\);
    
    un1_state_39_1_0_a3_0_1 : CFG3
      generic map(INIT => x"10")

      port map(A => \ins1[25]_net_1\, B => \ins1[24]_net_1\, C
         => \state[25]_net_1\, Y => \un1_state_39_1_0_a3_0_1\);
    
    \mask[4]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(4), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[4]_net_1\);
    
    \d_HADDR_0_iv_0_0_0[24]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_22_S, B => 
        \d_HADDR_0_iv_0_0_a3_0_0[24]_net_1\, C => HREADY_i_3, D
         => un1_state_30, Y => \d_HADDR_0_iv_0_0_0[24]_net_1\);
    
    \ins1[26]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(26), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[26]_net_1\);
    
    \count_RNI0JMT[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_266, B => \count[1]_net_1\, Y => 
        \d_count_0_a3_3_0[1]\);
    
    \state[13]\ : SLE
      port map(D => \state[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        HREADY_i_3_i_0, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[13]_net_1\);
    
    \expected[7]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(7), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[7]_net_1\);
    
    \haddr_write[3]\ : SLE
      port map(D => un46_d_haddr_cry_3_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[3]_net_1\);
    
    \count_RNI5T641[0]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => N_2570, B => \count[0]_net_1\, C => N_317, D
         => N_249, Y => N_2061);
    
    \HWDATA_int_RNO_1[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \state[10]_net_1\, B => \acc[20]_net_1\, Y
         => N_485);
    
    \or_br.d_busy\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \envm_soft_reset[1]_net_1\, B => 
        \envm_soft_reset[0]_net_1\, C => \envm_busy[1]_net_1\, D
         => \envm_busy[0]_net_1\, Y => d_busy);
    
    \HWDATA_int_RNO_1[25]\ : CFG4
      generic map(INIT => x"8A00")

      port map(A => d_HWDATA_0_iv_5_1424_a8_0_0, B => 
        \count[0]_net_1\, C => N_249, D => N_251, Y => N_2400);
    
    \mask[14]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(14), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[14]_net_1\);
    
    \state_RNIVVQK[22]\ : CFG2
      generic map(INIT => x"8")

      port map(A => d_state_1_sqmuxa_1_i_0, B => 
        \state[22]_net_1\, Y => N_4687);
    
    \d_acc_0[20]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[20]_net_1\, B => \ins2[20]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(20), D => \state[8]_net_1\, Y => 
        N_1157);
    
    \haddr_fetch_RNO[11]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_9_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[11]\, D => N_4812, Y => N_119_i_0);
    
    \rdata_RNI74OE[31]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \state[22]_net_1\, B => \rdata[31]_net_1\, Y
         => d_HWDATA_0_iv_1640_a8_3_0);
    
    \state[15]\ : SLE
      port map(D => \state_ns[13]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[15]_net_1\);
    
    \state[18]\ : SLE
      port map(D => \state[19]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        HREADY_i_3_i_0, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[18]_net_1\);
    
    \count[1]\ : SLE
      port map(D => \d_count[1]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[1]_net_1\);
    
    \rdata[15]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(15), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[15]_net_1\);
    
    \HADDR_int[30]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[30]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[30]\);
    
    d_HWRITE_0_sqmuxa_4_0_a3 : CFG2
      generic map(INIT => x"4")

      port map(A => \bytecount[0]_net_1\, B => 
        \bytecount[1]_net_1\, Y => N_661);
    
    \pause_count_RNO[3]\ : CFG4
      generic map(INIT => x"00AD")

      port map(A => \pause_count[3]_net_1\, B => 
        \pause_count[4]_net_1\, C => N_4811, D => N_3400, Y => 
        N_4808_i_0);
    
    \d_HADDR_0_iv_2[4]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[4]_net_1\, B => \ins2[4]_net_1\, 
        C => N_4873, D => N_4874, Y => \d_HADDR_0_iv_2[4]_net_1\);
    
    \bytecount[8]\ : SLE
      port map(D => N_42_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[8]_net_1\);
    
    \ins1[7]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(7), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[7]_net_1\);
    
    \haddr_fetch[15]\ : SLE
      port map(D => N_4342_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[15]_net_1\);
    
    \d_acc_1[5]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[5]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(5), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[5]\);
    
    \d_acc[14]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1151, C => 
        \ins2[14]_net_1\, D => \acc[14]_net_1\, Y => 
        \d_acc[14]_net_1\);
    
    \rdata[12]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(12), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[12]_net_1\);
    
    \haddr_fetch_RNO[19]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_17_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[19]\, D => N_4812, Y => 
        N_4367_i_0);
    
    \haddr_fetch_RNO[16]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_14_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[16]\, D => N_4812, Y => 
        N_4719_i_0);
    
    opcode_0_a3_0_0_a2 : CFG3
      generic map(INIT => x"01")

      port map(A => \ins1[26]_net_1\, B => \ins1[24]_net_1\, C
         => N_80, Y => N_198);
    
    d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0 : CFG2
      generic map(INIT => x"2")

      port map(A => \bytecount[0]_net_1\, B => 
        \bytecount[1]_net_1\, Y => 
        \d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0\);
    
    \acc[28]\ : SLE
      port map(D => \d_acc[28]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[28]_net_1\);
    
    un1_state_30_0_o3 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \state[26]_net_1\, B => \ins1[31]_net_1\, C
         => \state[21]_net_1\, D => N_109_i, Y => N_4814);
    
    \count_RNO_1[1]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => \d_count_0_0_0[1]\, B => N_319, C => N_375, D
         => \d_count_0_a2_1_c_1[1]\, Y => \d_count_0_2[1]\);
    
    \mask[22]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(22), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[22]_net_1\);
    
    un46_d_haddr_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \HADDR_int_fast[0]_net_1\, B => 
        \ins1[16]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        GND_net_1, S => OPEN, Y => un46_d_haddr_cry_0_Y, FCO => 
        \un46_d_haddr_cry_0\);
    
    \count_RNO_3[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => N_444, B => \d_count_0_0_tz[1]\, C => N_109_i, 
        Y => \d_count_0_0_0[1]\);
    
    \d_HADDR_0_iv_2[9]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_9_S, B => 
        \d_HADDR_0_iv_0[9]_net_1\, C => \ins2_m[9]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[9]_net_1\);
    
    un46_d_haddr_cry_30_1 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[7]\, B => 
        \ConfigMaster_0_M_HADDR[4]\, C => 
        \ConfigMaster_0_M_HADDR[5]\, D => 
        \ConfigMaster_0_M_HADDR[6]\, FCI => 
        un46_d_haddr_cry_3_0_FCO, S => OPEN, Y => OPEN, FCO => 
        un46_d_haddr_cry_30_1_FCO);
    
    \rdata[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[1]_net_1\);
    
    un46_d_haddr_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[15]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_14\, S => un46_d_haddr_s_15_S, Y => 
        OPEN, FCO => OPEN);
    
    un1_rdata_0_I_57 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[13]_net_1\, B => N_343_i, C => 
        \expected[13]_net_1\, D => \mask[13]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[5]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[6]\);
    
    \ins1[30]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(30), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[30]_net_1\);
    
    \d_ins2[12]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(12), B => un28_opcode, 
        Y => \d_ins2[12]_net_1\);
    
    \acc[10]\ : SLE
      port map(D => \d_acc[10]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[10]_net_1\);
    
    un1_rdata_0_I_87 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[3]_net_1\, B => N_347_i, C => 
        \expected[3]_net_1\, D => \mask[3]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[0]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[1]\);
    
    \d_HADDR_0_iv_1[11]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_0[11]_net_1\, B => 
        \haddr_fetch[11]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1[11]_net_1\);
    
    \bytecount_RNO[4]\ : CFG3
      generic map(INIT => x"70")

      port map(A => \state[21]_net_1\, B => N_109_i, C => N_105, 
        Y => N_34_i_0);
    
    un7_hready_2_RNIHUMF1 : CFG2
      generic map(INIT => x"E")

      port map(A => N_4777_1, B => N_403, Y => N_277);
    
    \haddr_write[27]\ : SLE
      port map(D => un46_d_haddr_cry_27_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[27]_net_1\);
    
    \count_RNO_1[0]\ : CFG4
      generic map(INIT => x"BE00")

      port map(A => \d_count_i_a2_2_1_0[0]\, B => 
        \count[0]_net_1\, C => HREADY_i_3, D => 
        \d_count_i_a2_2_1[0]\, Y => N_452);
    
    \haddr_write[10]\ : SLE
      port map(D => un46_d_haddr_cry_10_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[10]_net_1\);
    
    \ins2[16]\ : SLE
      port map(D => \d_ins2[16]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[16]_net_1\);
    
    un13_d_haddr_1_cry_16 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[18]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_15\, S => un13_d_haddr_1_cry_16_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_16\);
    
    \state_RNO[24]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \state[24]_net_1\, B => N_78, C => HREADY_i_3, 
        Y => N_12_i_0);
    
    \state_ns_0_rep1[7]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \state_21_rep1\, B => d_state_1_sqmuxa_1_i_0, 
        C => N_109_i, D => N_101, Y => \state_ns_rep1[7]\);
    
    \expected[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[1]_net_1\);
    
    \bytecount_RNO[12]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_114, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_50_i_0);
    
    \d_HADDR_0_iv_0_fast[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[0]_net_1\, C => \haddr_fetch[0]_net_1\, 
        Y => \d_HADDR_fast[0]\);
    
    \haddr_fetch_RNO[4]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_2_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[4]\, D => N_4812, Y => N_2921_i_0);
    
    \envm_busy[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_14_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \envm_busy[0]_net_1\);
    
    \state_RNI9A211[22]\ : CFG3
      generic map(INIT => x"5D")

      port map(A => N_274, B => N_251, C => N_249, Y => N_258);
    
    un1_d_HWRITE_0_sqmuxa_0_1 : CFG4
      generic map(INIT => x"0001")

      port map(A => \bytecount[3]_net_1\, B => 
        \d_HTRANS_0_sqmuxa_4_1_1_o3_1\, C => \bytecount[5]_net_1\, 
        D => \bytecount[4]_net_1\, Y => 
        \un1_d_HWRITE_0_sqmuxa_0_1\);
    
    \un7_iv_0_a1_0_RNIS4RTN[14]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un7_iv_0_a1_0[14]_net_1\, B => 
        \count[1]_net_1\, C => d_m2_e_1, D => 
        defSlaveSMNextState_m_0_3, Y => N_541);
    
    un1_state_46_0 : CFG4
      generic map(INIT => x"ECCC")

      port map(A => \ins1[31]_net_1\, B => \state[15]_net_1\, C
         => \un1_d_HWRITE_0_sqmuxa\, D => \state[22]_net_1\, Y
         => \un1_state_46_0\);
    
    \state_ns_i_0_o2_0[21]\ : CFG4
      generic map(INIT => x"005B")

      port map(A => \ins1[26]_net_1\, B => \ins1[24]_net_1\, C
         => \ins1[25]_net_1\, D => N_80, Y => N_379);
    
    \state_ns_0[11]\ : CFG4
      generic map(INIT => x"FCFA")

      port map(A => \state[18]_net_1\, B => \state[17]_net_1\, C
         => \state[15]_net_1\, D => HREADY_i_3, Y => 
        \state_ns[11]\);
    
    \state_ns_i_0_x2_1[1]\ : CFG4
      generic map(INIT => x"FFE4")

      port map(A => \ins1[26]_net_1\, B => \ins1[24]_net_1\, C
         => \ins1[25]_net_1\, D => N_80, Y => N_93_i);
    
    \count_RNIDU2E[0]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \state[21]_net_1\, B => N_249, C => 
        \count[0]_net_1\, Y => N_656);
    
    \d_HADDR_0_iv[27]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \un13_d_haddr_1_m[27]\, B => 
        un46_d_haddr_cry_27_S, C => \d_HADDR_0_iv_1_0[27]_net_1\, 
        D => N_247, Y => \d_HADDR[27]\);
    
    \acc[19]\ : SLE
      port map(D => \d_acc[19]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[19]_net_1\);
    
    \envm_soft_reset[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_696_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \envm_soft_reset[1]_net_1\);
    
    \state_ns_i_0_a2_3_0_1[1]\ : CFG4
      generic map(INIT => x"22F2")

      port map(A => N_917, B => N_156, C => N_117, D => 
        \state_ns_i_a2_10_i_2[1]_net_1\, Y => 
        \state_ns_i_0_a2_3_0_1[1]_net_1\);
    
    \haddr_fetch_RNO[9]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_7_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[9]\, D => N_4812, Y => N_4418_i_0);
    
    \count_RNI7TNO3[0]\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => d_HWDATA_0_iv_25_605_7_1_1, B => N_47, C => 
        \count[0]_net_1\, D => N_249, Y => N_2246_1);
    
    \HWDATA_int_RNO[5]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_25_605_7_1, B => N_2246_1, C
         => \rdata[5]_net_1\, D => N_403, Y => 
        \HWDATA_int_RNO[5]_net_1\);
    
    \state_RNO[14]\ : CFG4
      generic map(INIT => x"AA0C")

      port map(A => \state[14]_net_1\, B => N_191, C => N_198, D
         => HREADY_i_3, Y => N_16_i_0);
    
    \state_RNIP2C0P[22]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => HREADY_i_3, B => \d_count_0_o3_3_1[1]\, C => 
        N_251, Y => N_375);
    
    \count_RNO_0[0]\ : CFG3
      generic map(INIT => x"02")

      port map(A => N_259, B => N_251, C => HREADY_i_3, Y => 
        N_453);
    
    \HWDATA_int_RNO[18]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_12_1118_0_0, B => N_286, C => 
        \rdata[18]_net_1\, D => N_283, Y => 
        \HWDATA_int_RNO[18]_net_1\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_a2_0_RNO : CFG4
      generic map(INIT => x"0048")

      port map(A => \count[0]_net_1\, B => \state[21]_net_1\, C
         => \count[1]_net_1\, D => defSlaveSMNextState_m_0_2, Y
         => un1_m3_e_1);
    
    \HADDR_int[6]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[6]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[6]\);
    
    \haddr_fetch_RNO[6]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_4_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[6]\, D => N_4812, Y => N_4720_i_0);
    
    \d_HADDR_0_iv_0_2_RNO[17]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \ins2[17]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_i_m[17]\);
    
    \d_HADDR_0_iv_2[2]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_2_S, B => 
        \d_HADDR_0_iv_0[2]_net_1\, C => \ins2_m[2]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[2]_net_1\);
    
    \d_HADDR_0_iv_0[7]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_0_1[7]_net_1\, B => 
        un46_d_haddr_cry_7_S, C => \d_HADDR_0_iv_0_1_0[7]_net_1\, 
        D => N_247, Y => \d_HADDR[7]\);
    
    \d_HADDR_0_iv_2_RNO[19]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[19]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[19]\);
    
    \state_ns_0[2]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \state[26]_net_1\, B => \state[27]_net_1\, C
         => N_929, D => HREADY_i_3, Y => \state_ns[2]\);
    
    \expected[6]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(6), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[6]_net_1\);
    
    un13_d_haddr_1_s_29 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[31]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_28\, S => un13_d_haddr_1_s_29_S, Y
         => OPEN, FCO => OPEN);
    
    \ins1[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[1]_net_1\);
    
    \mask[11]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(11), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[11]_net_1\);
    
    \haddr_fetch_RNO[13]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_11_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[13]\, D => N_4812, Y => 
        \haddr_fetch_RNO[13]_net_1\);
    
    \HWDATA_int_RNO[28]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => d_HWDATA_0_iv_2_1532_5_0, B => 
        \rdata[28]_net_1\, C => N_686_2, D => N_277, Y => 
        \HWDATA_int_RNO[28]_net_1\);
    
    un13_d_haddr_1_cry_24 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[26]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_23\, S => un13_d_haddr_1_cry_24_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_24\);
    
    \state_ns_0_o2[8]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \state[12]_net_1\, B => \state[9]_net_1\, C
         => N_138, D => N_789, Y => N_133);
    
    un13_d_haddr_1_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[14]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_11\, S => un13_d_haddr_1_s_12_S, Y
         => OPEN, FCO => OPEN);
    
    \d_ins2[31]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(31), B => un28_opcode, 
        Y => \d_ins2[31]_net_1\);
    
    \acc[25]\ : SLE
      port map(D => \d_acc[25]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[25]_net_1\);
    
    \haddr_fetch[18]\ : SLE
      port map(D => \haddr_fetch_RNO[18]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[18]_net_1\);
    
    \rdata[11]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(11), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[11]_net_1\);
    
    \state_RNI7N251[22]\ : CFG4
      generic map(INIT => x"50DC")

      port map(A => N_274, B => N_251, C => N_252, D => N_249, Y
         => N_255);
    
    \rdata[24]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(24), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[24]_net_1\);
    
    \bytecount[9]\ : SLE
      port map(D => N_44_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[9]_net_1\);
    
    \d_ins2[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(2), B => un28_opcode, 
        Y => \d_ins2[2]_net_1\);
    
    \state[5]\ : SLE
      port map(D => \state[6]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[5]_net_1\);
    
    \state[20]\ : SLE
      port map(D => \state_ns[8]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[20]_net_1\);
    
    \mask[29]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(29), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[29]_net_1\);
    
    \acc[26]\ : SLE
      port map(D => \d_acc[26]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[26]_net_1\);
    
    \HADDR_int[2]\ : SLE
      port map(D => \d_HADDR[2]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[2]\);
    
    un1_rdata_0_I_52 : CFG3
      generic map(INIT => x"6A")

      port map(A => \expected[9]_net_1\, B => \rdata[9]_net_1\, C
         => \mask[9]_net_1\, Y => un1_rdata_0_N_37);
    
    d_HWDATA_0_sqmuxa_2_RNID7K81 : CFG4
      generic map(INIT => x"020E")

      port map(A => N_251, B => \state[10]_net_1\, C => 
        \d_HWDATA_0_sqmuxa_2\, D => HREADY_i_3, Y => 
        un1_state_38_i_0);
    
    \HWDATA_int[6]\ : SLE
      port map(D => \HWDATA_int_RNO[6]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(6));
    
    \rdata[23]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(23), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[23]_net_1\);
    
    \rdata[30]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(30), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[30]_net_1\);
    
    \state_RNIHO0QN[23]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => defSlaveSMNextState_m_0_2, B => 
        \state[23]_net_1\, C => un1_state_31_i_i_a2_0_d_1_0_1, D
         => defSlaveSMNextState_m_0_3, Y => N_4874);
    
    \HADDR_int[22]\ : SLE
      port map(D => \d_HADDR[22]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[22]\);
    
    un1_rdata_0_I_82 : CFG3
      generic map(INIT => x"6A")

      port map(A => \expected[5]_net_1\, B => \rdata[5]_net_1\, C
         => \mask[5]_net_1\, Y => un1_rdata_0_N_12);
    
    state_m2_e_1 : CFG4
      generic map(INIT => x"A0A8")

      port map(A => \state_m2_e_0\, B => N_117, C => N_917, D => 
        \state_ns_i_a2_10_i_2[1]_net_1\, Y => \state_m2_e_1\);
    
    un13_d_haddr_1_cry_22 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[24]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_21\, S => un13_d_haddr_1_cry_22_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_22\);
    
    state_m3_i_a3 : CFG4
      generic map(INIT => x"040C")

      port map(A => \state_ns_i_0_a2_3_d_0[1]_net_1\, B => N_74, 
        C => N_198, D => \state_m2_e_2\, Y => \state_m3_i_a3\);
    
    \HWDATA_int_RNO[19]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_11_1163_0_0, B => N_288, C => 
        \rdata[19]_net_1\, D => N_283, Y => 
        \HWDATA_int_RNO[19]_net_1\);
    
    \d_HADDR_0_iv_0[9]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_7_S, B => 
        \haddr_write[9]_net_1\, C => N_4874, D => un1_state_30, Y
         => \d_HADDR_0_iv_0[9]_net_1\);
    
    \d_ins2[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(6), B => un28_opcode, 
        Y => \d_ins2[6]_net_1\);
    
    \HWDATA_int[22]\ : SLE
      port map(D => \HWDATA_int_RNO[22]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(22));
    
    \d_HADDR_0_iv_0_1[7]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[7]_net_1\, B => \ins2[7]_net_1\, 
        C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_0_1[7]_net_1\);
    
    \d_HADDR_0_iv_0_2[12]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_12_S, B => 
        \d_HADDR_0_iv_0_0[12]_net_1\, C => N_4445, D => N_247, Y
         => \d_HADDR_0_iv_0_2[12]_net_1\);
    
    \count_RNIHUMF1[1]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \count[1]_net_1\, B => N_403, C => N_262, Y
         => N_264);
    
    \HWDATA_int_RNO[29]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \acc[29]_net_1\, B => \state[10]_net_1\, C
         => N_301, D => d_HWDATA_0_iv_1_1568_0_1, Y => 
        \HWDATA_int_RNO[29]_net_1\);
    
    \d_HADDR_0_iv_0_0[3]\ : CFG4
      generic map(INIT => x"DDDC")

      port map(A => un13_d_haddr_1_cry_1_S, B => \state_ns[0]\, C
         => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0_0[3]_net_1\);
    
    \ins1_RNIUC04[22]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \ins1[23]_net_1\, B => \ins1[22]_net_1\, C
         => \ins1[21]_net_1\, D => \ins1[20]_net_1\, Y => N_252);
    
    \ins2[22]\ : SLE
      port map(D => \d_ins2[22]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[22]_net_1\);
    
    \acc[4]\ : SLE
      port map(D => \d_acc[4]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[4]_net_1\);
    
    \haddr_fetch[29]\ : SLE
      port map(D => N_18_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[29]_net_1\);
    
    \bytecount_RNO[13]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4341, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_52_i_0);
    
    \mask[10]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(10), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[10]_net_1\);
    
    \ins1[15]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(15), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[15]_net_1\);
    
    \d_HADDR_0_iv[29]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \un13_d_haddr_1_m[29]\, B => 
        un46_d_haddr_cry_29_S, C => \d_HADDR_0_iv_1_0[29]_net_1\, 
        D => N_247, Y => \d_HADDR[29]\);
    
    \ins1_RNIHBC1J1[2]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[2]_net_1\, B => N_78, C => N_164, 
        D => \ins1[2]_net_1\, FCI => d_bytecount_i_m2_cry_1, S
         => N_104, Y => OPEN, FCO => d_bytecount_i_m2_cry_2);
    
    un13_d_haddr_1_cry_21 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[23]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_20\, S => un13_d_haddr_1_cry_21_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_21\);
    
    \d_HADDR_0_iv_2[14]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[14]_net_1\, B => 
        \ins2[14]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_2[14]_net_1\);
    
    \acc[21]\ : SLE
      port map(D => \d_acc[21]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[21]_net_1\);
    
    \ins1[8]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(8), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[8]_net_1\);
    
    un13_d_haddr_1_cry_20 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[22]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_19\, S => un13_d_haddr_1_cry_20_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_20\);
    
    un46_d_haddr_cry_30_5 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[15]\, B => 
        \ConfigMaster_0_M_HADDR[12]\, C => 
        \ConfigMaster_0_M_HADDR[13]\, D => 
        \ConfigMaster_0_M_HADDR[14]\, FCI => 
        un46_d_haddr_cry_30_3_FCO, S => OPEN, Y => OPEN, FCO => 
        un46_d_haddr_cry_30_5_FCO);
    
    un1_rdata_0_I_44_i_0_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[18]_net_1\, B => \rdata[18]_net_1\, 
        C => \mask[18]_net_1\, Y => N_335_i);
    
    un1_d_HWRITE_1_sqmuxa_2_i_a2_0 : CFG4
      generic map(INIT => x"F0D0")

      port map(A => un1_m3_e_1, B => 
        un1_state_31_i_i_a2_0_d_1_0_1, C => 
        \un1_d_HWRITE_1_sqmuxa_2_i_a2_0_0\, D => 
        defSlaveSMNextState_m_0_3, Y => N_4901);
    
    \HADDR_int[11]\ : SLE
      port map(D => \d_HADDR[11]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[11]\);
    
    un1_rdata_0_I_8_i_x2_0 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[0]_net_1\, B => \rdata[0]_net_1\, C
         => \mask[0]_net_1\, Y => N_83_i);
    
    \d_HADDR_0_iv_1_1[31]\ : CFG3
      generic map(INIT => x"5D")

      port map(A => \d_HADDR_0_iv_1_0[31]_net_1\, B => 
        un46_d_haddr_s_31_S, C => N_247, Y => 
        \d_HADDR_0_iv_1_1[31]_net_1\);
    
    \d_ins2[22]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(22), B => un28_opcode, 
        Y => \d_ins2[22]_net_1\);
    
    \ins2[24]\ : SLE
      port map(D => \d_ins2[24]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[24]_net_1\);
    
    \HWDATA_int_RNO_1[17]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \state[10]_net_1\, B => \acc[17]_net_1\, Y
         => N_475);
    
    un1_hready_2_0 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => N_4912, B => N_252, C => 
        defSlaveSMNextState_m, D => un1_state_31_i_i_a2_0_d_1_0_1, 
        Y => un1_hready_2);
    
    \un1_d_state_1_sqmuxa_1_0_m2[0]\ : CFG4
      generic map(INIT => x"CCE4")

      port map(A => d_N_3_mux_0, B => d_state_1_sqmuxa_1_i_0, C
         => \ins1[31]_net_1\, D => N_266, Y => 
        \un1_d_state_1_sqmuxa_1[0]\);
    
    \haddr_fetch[16]\ : SLE
      port map(D => N_4719_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[16]_net_1\);
    
    \d_ins2[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(15), B => un28_opcode, 
        Y => \d_ins2[15]_net_1\);
    
    \d_ins2[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(4), B => un28_opcode, 
        Y => \d_ins2[4]_net_1\);
    
    \d_HADDR_0_iv_0_2[30]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => \haddr_write[30]_net_1\, B => 
        \ins2[30]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_0_2[30]_net_1\);
    
    un1_rdata_0_I_35 : CFG3
      generic map(INIT => x"6A")

      port map(A => \expected[20]_net_1\, B => \rdata[20]_net_1\, 
        C => \mask[20]_net_1\, Y => un1_rdata_0_N_53);
    
    \HWDATA_int_RNO_0[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[8]_net_1\, D => \rdata[24]_net_1\, Y => 
        d_HWDATA_0_iv_22_740_6_0);
    
    \count_RNO_9[0]\ : CFG4
      generic map(INIT => x"2033")

      port map(A => \state[21]_net_1\, B => \count[0]_net_1\, C
         => N_109_i, D => N_542_2, Y => \d_count_i_0[0]\);
    
    \state_ns_0_0[17]\ : CFG4
      generic map(INIT => x"D5C0")

      port map(A => \ins1[24]_net_1\, B => \state[11]_net_1\, C
         => HREADY_i_3, D => N_411_2, Y => \state_ns[17]\);
    
    \count_RNIOOC0O[0]\ : CFG4
      generic map(INIT => x"0DDD")

      port map(A => \d_count_0_a3_8_0[1]\, B => \count[0]_net_1\, 
        C => d_m2_e_1, D => d_m2_e_2_0_1, Y => d_m2_e_2_0);
    
    \d_HADDR_0_iv_2_RNO[28]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[28]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[28]\);
    
    \HWDATA_int[31]\ : SLE
      port map(D => \HWDATA_int_RNO[31]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(31));
    
    state_m3_i_8 : CFG4
      generic map(INIT => x"EAEE")

      port map(A => \state_m3_i_7\, B => HREADY_i_3, C => 
        \state[25]_net_1\, D => N_917, Y => \state_m3_i_8\);
    
    \rdata_RNIF5VS1[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[20]_net_1\, B => \rdata[4]_net_1\, C
         => N_592, D => N_254, Y => N_686_2);
    
    un46_d_haddr_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[18]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[2]\, C => GND_net_1, D => 
        GND_net_1, FCI => \un46_d_haddr_cry_1\, S => 
        un46_d_haddr_cry_2_S, Y => OPEN, FCO => 
        \un46_d_haddr_cry_2\);
    
    \d_HADDR_0_iv[28]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[28]_net_1\, C => \haddr_fetch[28]_net_1\, 
        Y => \d_HADDR[28]\);
    
    \ins2[4]\ : SLE
      port map(D => \d_ins2[4]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[4]_net_1\);
    
    d_count_1_sqmuxa_i_a2_0_o2_i_o2_RNIPVPC4 : CFG4
      generic map(INIT => x"20A0")

      port map(A => d_N_3_mux_0, B => N_281, C => N_259, D => 
        \d_count_0_a3_3_0[1]\, Y => \d_count_0_a2_1_2_1[1]\);
    
    un1_d_HWRITE_0_sqmuxa_2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_d_HWRITE_0_sqmuxa_2_0_0\, B => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => un1_d_HWRITE_0_sqmuxa_2);
    
    \d_ins2[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(7), B => un28_opcode, 
        Y => \d_ins2[7]_net_1\);
    
    \ins2[0]\ : SLE
      port map(D => \d_ins2[0]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[0]_net_1\);
    
    un46_d_haddr_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[14]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_13\, S => un46_d_haddr_cry_14_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_14\);
    
    \d_acc_1[10]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[10]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(10), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[10]\);
    
    un1_hready_2_0_0 : CFG3
      generic map(INIT => x"FD")

      port map(A => N_252, B => un1_state_31_i_i_a2_0_d_1_0_1, C
         => N_4912, Y => \un1_hready_2_0_0\);
    
    \state_RNIN40R[22]\ : CFG4
      generic map(INIT => x"EC00")

      port map(A => \state[22]_net_1\, B => \state[21]_net_1\, C
         => N_252, D => N_249, Y => N_257);
    
    \HWDATA_int[30]\ : SLE
      port map(D => N_2525, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(30));
    
    \d_acc[22]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1159, C => 
        \ins2[22]_net_1\, D => \acc[22]_net_1\, Y => 
        \d_acc[22]_net_1\);
    
    \state_ns_0_a2_0_1[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \state[21]_net_1\, B => 
        d_state_1_sqmuxa_1_i_0, C => N_109_i, Y => 
        \state_ns_0_a2_0_1[5]_net_1\);
    
    \HWDATA_int[25]\ : SLE
      port map(D => \HWDATA_int_RNO[25]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(25));
    
    \d_HADDR_0_iv_0[10]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[10]_net_1\, C => 
        \haddr_fetch[10]_net_1\, Y => \d_HADDR[10]\);
    
    \ins2[6]\ : SLE
      port map(D => \d_ins2[6]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[6]_net_1\);
    
    un28_opcode_0 : CFG4
      generic map(INIT => x"007B")

      port map(A => \ins1[26]_net_1\, B => \ins1[24]_net_1\, C
         => \ins1[25]_net_1\, D => N_80, Y => un28_opcode);
    
    \HADDR_int[29]\ : SLE
      port map(D => \d_HADDR[29]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[29]\);
    
    \count_RNID2MUO[0]\ : CFG4
      generic map(INIT => x"084C")

      port map(A => HREADY_i_3, B => d_m2_e_2_0, C => 
        \d_count_0_a3_8_0[1]\, D => N_591, Y => d_m2_e_2_2);
    
    \expected[12]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(12), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[12]_net_1\);
    
    \rdata[16]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(16), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[16]_net_1\);
    
    \ins1_RNIU9N0C2[3]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[3]_net_1\, B => N_78, C => N_164, 
        D => \ins1[3]_net_1\, FCI => d_bytecount_i_m2_cry_2, S
         => N_1104, Y => OPEN, FCO => d_bytecount_i_m2_cry_3);
    
    \state_ns_a2_i_i_a2[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => \state[17]_net_1\, Y => 
        N_480);
    
    \HWDATA_int_RNO_2[30]\ : CFG3
      generic map(INIT => x"37")

      port map(A => N_4777_1, B => \rdata[30]_net_1\, C => N_403, 
        Y => d_HWDATA_0_iv_0_1604_1_0);
    
    un13_d_haddr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[16]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_13\, S => un13_d_haddr_1_cry_14_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_14\);
    
    \d_HADDR_0_iv[20]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[20]_net_1\, C => \haddr_fetch[20]_net_1\, 
        Y => \d_HADDR[20]\);
    
    un46_d_haddr_axb_0 : CFG2
      generic map(INIT => x"6")

      port map(A => \HADDR_int_fast[0]_net_1\, B => 
        \ins1[16]_net_1\, Y => \un46_d_haddr_axb_0\);
    
    pause_count_n3_i_o2_RNIKOEU : CFG3
      generic map(INIT => x"F7")

      port map(A => \pause_count[4]_net_1\, B => 
        \pause_count[3]_net_1\, C => N_4811, Y => N_4813);
    
    \mask[8]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(8), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[8]_net_1\);
    
    un1_rdata_0_I_62_i_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[12]_net_1\, B => \rdata[12]_net_1\, 
        C => \mask[12]_net_1\, Y => N_343_i);
    
    \d_HADDR_0_iv_0_0[21]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_19_S, B => 
        \haddr_write[21]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[21]_net_1\);
    
    \ins1_RNIHHOUM4[6]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[6]_net_1\, B => N_78, C => N_164, 
        D => \ins1[6]_net_1\, FCI => d_bytecount_i_m2_cry_5, S
         => N_4336, Y => OPEN, FCO => d_bytecount_i_m2_cry_6);
    
    \ins1[4]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(4), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[4]_net_1\);
    
    \d_ins2[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(8), B => un28_opcode, 
        Y => \d_ins2[8]_net_1\);
    
    \state_ns_0_0[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \ins1[24]_net_1\, B => \state[8]_net_1\, C
         => HREADY_i_3, D => N_411_2, Y => \state_ns[20]\);
    
    un46_d_haddr_cry_26 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[26]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_25\, S => un46_d_haddr_cry_26_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_26\);
    
    un1_state_42_0_a3_1_1 : CFG4
      generic map(INIT => x"0004")

      port map(A => defSlaveSMNextState_m_0_2, B => N_117, C => 
        un1_state_31_i_i_a2_0_d_1_0_1, D => 
        defSlaveSMNextState_m_0_3, Y => N_182_1);
    
    \state_ns_a2_1_i_o2[4]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_93_i, B => N_86, Y => N_96);
    
    \ins1[22]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(22), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[22]_net_1\);
    
    \d_acc_1_0[4]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[4]_net_1\, B => \acc[4]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[4]_net_1\);
    
    \haddr_write[5]\ : SLE
      port map(D => un46_d_haddr_cry_5_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[5]_net_1\);
    
    un13_d_haddr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[7]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_4\, S => un13_d_haddr_1_cry_5_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_5\);
    
    \d_acc_0[9]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[9]_net_1\, B => \ins2[9]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(9), D => \state[8]_net_1\, Y => 
        N_1146);
    
    \HADDR_int_RNO[15]\ : CFG4
      generic map(INIT => x"5040")

      port map(A => \un13_d_haddr_1_i_m[15]\, B => 
        un46_d_haddr_s_15_S, C => \d_HADDR_0_iv_i_1[15]\, D => 
        N_247, Y => \d_HADDR_0_iv_i_0[15]\);
    
    \d_acc_0[25]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[25]_net_1\, B => \ins2[25]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(25), D => \state[8]_net_1\, Y => 
        N_1162);
    
    \HWDATA_int_RNO[1]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_29_425_0_0, B => N_296, C => 
        \rdata[17]_net_1\, D => N_271, Y => 
        \HWDATA_int_RNO[1]_net_1\);
    
    \count_RNO_3[0]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \count[0]_net_1\, B => N_369, C => HREADY_i_3, 
        Y => N_450);
    
    \haddr_write[22]\ : SLE
      port map(D => un46_d_haddr_cry_22_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[22]_net_1\);
    
    \d_acc_1[28]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_789, B => \d_acc_1_0[28]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(28), Y => \d_acc[28]\);
    
    \d_HADDR_0_iv[14]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_2[14]_net_1\, B => 
        un46_d_haddr_cry_14_S, C => \d_HADDR_0_iv_1[14]_net_1\, D
         => N_247, Y => \d_HADDR[14]\);
    
    \HWDATA_int_RNO_0[18]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_601, C => 
        \acc[18]_net_1\, D => \rdata[2]_net_1\, Y => 
        d_HWDATA_0_iv_12_1118_0_0);
    
    \acc[3]\ : SLE
      port map(D => \d_acc[3]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[3]_net_1\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o2_1 : CFG4
      generic map(INIT => x"7773")

      port map(A => \state[22]_net_1\, B => N_251, C => 
        defSlaveSMNextState_m, D => 
        un1_d_HWRITE_1_sqmuxa_2_i_o3_1_2, Y => 
        \un1_d_HWRITE_1_sqmuxa_2_i_o2_1\);
    
    \rdata_RNI81HO[13]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \rdata[29]_net_1\, B => \rdata[13]_net_1\, C
         => \count[1]_net_1\, D => N_317, Y => N_4525);
    
    \bytecount[4]\ : SLE
      port map(D => N_34_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[4]_net_1\);
    
    \d_HADDR_0_iv[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[9]_net_1\, C => \haddr_fetch[9]_net_1\, Y
         => \d_HADDR[9]\);
    
    \state_RNI8PP21[22]\ : CFG4
      generic map(INIT => x"40FF")

      port map(A => \count[1]_net_1\, B => \state[22]_net_1\, C
         => N_276, D => N_263, Y => N_278);
    
    \ins2[30]\ : SLE
      port map(D => \d_ins2[30]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[30]_net_1\);
    
    \haddr_write[15]\ : SLE
      port map(D => un46_d_haddr_s_15_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[15]_net_1\);
    
    \ins1_RNI6F12Q[1]\ : ARI1
      generic map(INIT => x"5E44E")

      port map(A => \bytecount[1]_net_1\, B => N_78, C => 
        \ins1[1]_net_1\, D => \un7_iv[14]_net_1\, FCI => 
        d_bytecount_i_m2_cry_0, S => N_1102, Y => OPEN, FCO => 
        d_bytecount_i_m2_cry_1);
    
    \haddr_write[6]\ : SLE
      port map(D => un46_d_haddr_cry_6_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[6]_net_1\);
    
    \haddr_write[0]\ : SLE
      port map(D => un46_d_haddr_cry_0_Y, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[0]_net_1\);
    
    \HWDATA_int_RNO_2[27]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[22]_net_1\, B => \rdata[11]_net_1\, C
         => N_276, D => \count[1]_net_1\, Y => N_4431);
    
    \acc[17]\ : SLE
      port map(D => \d_acc[17]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[17]_net_1\);
    
    \d_HADDR_0_iv_2[25]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_25_S, B => 
        \d_HADDR_0_iv_0[25]_net_1\, C => \ins2_m[25]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[25]_net_1\);
    
    un13_d_haddr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[13]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_10\, S => un13_d_haddr_1_cry_11_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_11\);
    
    \ins1[24]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(24), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[24]_net_1\);
    
    un46_d_haddr_cry_19 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[19]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_18\, S => un46_d_haddr_cry_19_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_19\);
    
    \HADDR_int_RNO_0[15]\ : CFG3
      generic map(INIT => x"54")

      port map(A => un13_d_haddr_1_cry_13_S, B => 
        \un1_state_30_0_0\, C => N_4814, Y => 
        \un13_d_haddr_1_i_m[15]\);
    
    \state_ns_0[24]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \state[5]_net_1\, B => \state[4]_net_1\, C
         => HREADY_i_3, Y => \state_ns[24]\);
    
    \rdata_RNIMR2M[14]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \rdata[14]_net_1\, B => \rdata[6]_net_1\, C
         => \count[1]_net_1\, D => N_249, Y => 
        d_HWDATA_0_iv_8_1298_1_o2_i_m2_ns_1);
    
    \count_RNI3765[0]\ : CFG3
      generic map(INIT => x"5D")

      port map(A => \count[1]_net_1\, B => N_249, C => 
        \count[0]_net_1\, Y => N_4879);
    
    un1_rdata_0_I_21 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[14]_net_1\, B => N_339_i, C => 
        \expected[14]_net_1\, D => \mask[14]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[6]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[7]\);
    
    \d_acc_0[17]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[17]_net_1\, B => \ins2[17]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(17), D => \state[8]_net_1\, Y => 
        N_1154);
    
    \state_ns_i_0_a2_3_0[1]\ : CFG4
      generic map(INIT => x"5FDF")

      port map(A => N_86, B => \state[25]_net_1\, C => 
        \state_ns_i_0_a2_3_0_1[1]_net_1\, D => N_93_i, Y => N_74);
    
    \haddr_fetch_RNO[31]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_s_29_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[31]\, D => N_4812, Y => 
        N_4366_i_0);
    
    un13_d_haddr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[12]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_9\, S => un13_d_haddr_1_cry_10_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_10\);
    
    \haddr_write[8]\ : SLE
      port map(D => un46_d_haddr_cry_8_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[8]_net_1\);
    
    \haddr_fetch_RNO[3]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_1_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[3]\, D => N_4812, Y => N_53_i_0);
    
    \d_HADDR_0_iv_1[22]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[22]_net_1\, B => 
        \ins2[22]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_1[22]_net_1\);
    
    \ins1[11]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(11), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[11]_net_1\);
    
    \haddr_fetch_RNO[24]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_22_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[24]\, D => N_4812, Y => 
        \haddr_fetch_RNO[24]_net_1\);
    
    \d_acc_0[22]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[22]_net_1\, B => \ins2[22]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(22), D => \state[8]_net_1\, Y => 
        N_1159);
    
    d_HWRITE_0_sqmuxa_1_0_a3_1 : CFG3
      generic map(INIT => x"04")

      port map(A => \bytecount[2]_net_1\, B => N_661, C => N_249, 
        Y => \d_HWRITE_0_sqmuxa_1_0_a3_1\);
    
    \ins1[13]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(13), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[13]_net_1\);
    
    \HWDATA_int_RNO[3]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_27_515_0_0, B => N_288, C => 
        \rdata[19]_net_1\, D => N_271, Y => 
        \HWDATA_int_RNO[3]_net_1\);
    
    \state_ns_i_i_a3[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => N_259, Y => N_170);
    
    \d_acc_0[23]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[23]_net_1\, B => \ins2[23]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(23), D => \state[8]_net_1\, Y => 
        N_1160);
    
    \d_HADDR_0_iv_0[23]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_21_S, B => 
        \haddr_write[23]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[23]_net_1\);
    
    \d_HADDR_0_iv[25]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[25]_net_1\, C => \haddr_fetch[25]_net_1\, 
        Y => \d_HADDR[25]\);
    
    \ins1[18]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(18), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[18]_net_1\);
    
    \d_HADDR_0_iv_RNO[1]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \ConfigMaster_0_M_HADDR[1]\, B => 
        \un1_state_30_0_0\, C => N_4814, Y => 
        \un13_d_haddr_1_m[1]\);
    
    \d_HADDR_0_iv_2[8]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[8]_net_1\, B => \ins2[8]_net_1\, 
        C => N_4873, D => N_4874, Y => \d_HADDR_0_iv_2[8]_net_1\);
    
    \d_HADDR_0_iv_2_RNO[2]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[2]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[2]\);
    
    \d_HADDR_0_iv_0[5]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[5]_net_1\, C => \haddr_fetch[5]_net_1\, 
        Y => \d_HADDR[5]\);
    
    \count_RNIN95F1[1]\ : CFG4
      generic map(INIT => x"D0C0")

      port map(A => N_249, B => d_HWDATA_0_iv_20_812_o3_0_0, C
         => \count[1]_net_1\, D => N_251, Y => N_587);
    
    \state_ns_i_0_a2_3[1]\ : CFG4
      generic map(INIT => x"DD0D")

      port map(A => N_917, B => N_156, C => N_117, D => 
        \state_ns_i_a2_10_i_2[1]_net_1\, Y => N_148);
    
    \d_HADDR_0_iv_1[8]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_0[8]_net_1\, B => 
        \haddr_fetch[8]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1[8]_net_1\);
    
    \count_RNO_7[0]\ : CFG4
      generic map(INIT => x"CCCE")

      port map(A => N_674, B => \d_count_i_0[0]\, C => 
        \state[21]_net_1\, D => N_259, Y => \d_count_i_1[0]\);
    
    \acc[8]\ : SLE
      port map(D => \d_acc[8]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[8]_net_1\);
    
    \HWDATA_int_RNO[6]\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => d_HWDATA_0_iv_24_650_7_0, B => N_4891, C => 
        \rdata[22]_net_1\, D => N_4890, Y => 
        \HWDATA_int_RNO[6]_net_1\);
    
    d_mask_0_sqmuxa_i_i_a3 : CFG4
      generic map(INIT => x"0004")

      port map(A => defSlaveSMNextState_m_0_2, B => 
        \state[19]_net_1\, C => un1_state_31_i_i_a2_0_d_1_0_1, D
         => defSlaveSMNextState_m_0_3, Y => N_167);
    
    \d_HADDR_0_iv_0_0[18]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_16_S, B => 
        \haddr_write[18]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[18]_net_1\);
    
    \count_RNISU5S[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_257, B => N_585, Y => N_655);
    
    \HWDATA_int_RNO_1[21]\ : CFG4
      generic map(INIT => x"8F88")

      port map(A => \state[10]_net_1\, B => \acc[21]_net_1\, C
         => N_274, D => N_4541, Y => d_HWDATA_0_iv_9_1253_1_0);
    
    \d_ins2[25]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(25), B => un28_opcode, 
        Y => \d_ins2[25]_net_1\);
    
    \bytecount[15]\ : SLE
      port map(D => \d_bytecount[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[15]_net_1\);
    
    state_m2_e_2 : CFG4
      generic map(INIT => x"8CCC")

      port map(A => N_93_i, B => \state_m2_e_1\, C => 
        \state[25]_net_1\, D => N_97, Y => \state_m2_e_2\);
    
    \haddr_fetch[24]\ : SLE
      port map(D => \haddr_fetch_RNO[24]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[24]_net_1\);
    
    \HWDATA_int_RNO_1[27]\ : CFG4
      generic map(INIT => x"B3A0")

      port map(A => \state[10]_net_1\, B => N_263, C => 
        \acc[27]_net_1\, D => \rdata[11]_net_1\, Y => 
        d_HWDATA_0_iv_3_1496_0_0);
    
    \state[4]\ : SLE
      port map(D => \state_ns[24]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[4]_net_1\);
    
    \state_ns_0[9]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => N_4837, B => \state[19]_net_1\, C => 
        HREADY_i_3, Y => \state_ns[9]\);
    
    \d_HADDR_0_iv_0[8]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => un13_d_haddr_1_cry_6_S, B => \state[5]_net_1\, 
        C => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0[8]_net_1\);
    
    \ins2[12]\ : SLE
      port map(D => \d_ins2[12]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[12]_net_1\);
    
    \d_HADDR_0_iv_2[19]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_19_S, B => 
        \d_HADDR_0_iv_0[19]_net_1\, C => \ins2_m[19]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[19]_net_1\);
    
    \count_RNO[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \d_count_0_a2_1_d[1]\, B => \d_count_0_2[1]\, 
        C => N_445, Y => \d_count[1]\);
    
    \HADDR_int_RNO[6]\ : CFG4
      generic map(INIT => x"5040")

      port map(A => \d_HADDR_0_iv_2[6]_net_1\, B => 
        un46_d_haddr_cry_6_S, C => \d_HADDR_0_iv_i_1[6]\, D => 
        N_247, Y => \d_HADDR_0_iv_i_0[6]\);
    
    state_21_rep1_RNI4C9T : CFG4
      generic map(INIT => x"2A00")

      port map(A => \state_21_rep1\, B => masterDataInProg(0), C
         => CoreAHBLite_1_AHBmslave16_HREADY, D => 
        xhdl1328_i_m_0_1(0), Y => un1_state_31_i_i_a2_0_d_1_0_sx);
    
    \count_RNI5Q51[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \count[1]_net_1\, B => \count[0]_net_1\, Y
         => N_585);
    
    \d_HADDR_0_iv_2[20]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_20_S, B => 
        \d_HADDR_0_iv_0[20]_net_1\, C => \ins2_m[20]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[20]_net_1\);
    
    \rdata[2]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(2), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[2]_net_1\);
    
    \ins2[9]\ : SLE
      port map(D => \d_ins2[9]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[9]_net_1\);
    
    \haddr_fetch_RNO[20]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_18_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[20]\, D => N_4812, Y => 
        N_4560_i_0);
    
    \d_acc[15]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1152, C => 
        \ins2[15]_net_1\, D => \acc[15]_net_1\, Y => 
        \d_acc[15]_net_1\);
    
    un46_d_haddr_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[5]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_4\, S => un46_d_haddr_cry_5_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_5\);
    
    \HWDATA_int_RNO_0[16]\ : CFG4
      generic map(INIT => x"F8FF")

      port map(A => \acc[16]_net_1\, B => \state[10]_net_1\, C
         => N_4741, D => N_4889, Y => d_HWDATA_0_iv_14_1028_3_1);
    
    \rdata[18]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(18), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[18]_net_1\);
    
    \expected[22]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(22), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[22]_net_1\);
    
    \d_ins2[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(1), B => un28_opcode, 
        Y => \d_ins2[1]_net_1\);
    
    \count_RNIEROS[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => \count[1]_net_1\, B => N_4916, C => N_656, Y
         => N_254);
    
    un12_size_2_0_4 : CFG4
      generic map(INIT => x"0001")

      port map(A => \bytecount[15]_net_1\, B => 
        \bytecount[14]_net_1\, C => \bytecount[13]_net_1\, D => 
        \bytecount[12]_net_1\, Y => \un12_size_2_0_4\);
    
    \pause_count[4]\ : SLE
      port map(D => N_4809_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        pause_counte, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pause_count[4]_net_1\);
    
    un1_state_30_0_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \state[27]_net_1\, B => \state[25]_net_1\, C
         => \ins1[25]_net_1\, D => N_198, Y => \un1_state_30_0_0\);
    
    \ins1_RNIDA2053[4]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[4]_net_1\, B => N_78, C => N_164, 
        D => \ins1[4]_net_1\, FCI => d_bytecount_i_m2_cry_3, S
         => N_105, Y => OPEN, FCO => d_bytecount_i_m2_cry_4);
    
    \HADDR_int[12]\ : SLE
      port map(D => \d_HADDR[12]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[12]\);
    
    \ins2[14]\ : SLE
      port map(D => \d_ins2[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[14]_net_1\);
    
    \HWDATA_int[28]\ : SLE
      port map(D => \HWDATA_int_RNO[28]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(28));
    
    \rdata_RNIUQEJ1[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_4916, B => N_656, C => \rdata[17]_net_1\, D
         => N_388, Y => N_2380_3);
    
    un1_state_44_0_a3_1_RNISO1K : CFG4
      generic map(INIT => x"0001")

      port map(A => \un1_state_44_0_12\, B => N_4856, C => N_4854, 
        D => N_4857, Y => un1_state_44_i_0);
    
    un1_rdata_0_I_39 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[19]_net_1\, B => N_335_i, C => 
        \expected[19]_net_1\, D => \mask[19]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[8]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[9]\);
    
    \state[10]\ : SLE
      port map(D => \state[11]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        HREADY_i_3_i_0, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[10]_net_1\);
    
    \HWDATA_int_RNO_0[2]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_270, C => 
        \acc[2]_net_1\, D => \rdata[2]_net_1\, Y => 
        d_HWDATA_0_iv_28_470_3_0);
    
    \bytecount_RNO[14]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_116, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_55_i_0);
    
    \haddr_fetch[13]\ : SLE
      port map(D => \haddr_fetch_RNO[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[13]_net_1\);
    
    \mask[1]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(1), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[1]_net_1\);
    
    un1_state_39 : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \state[21]_net_1\, B => N_191, C => 
        \un1_state_39_1\, D => \un1_d_state_1_sqmuxa_1[0]\, Y => 
        \un1_state_39\);
    
    \d_acc_1_0[24]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_789, B => \d_acc_1_0_0[24]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(24), Y => \d_acc[24]\);
    
    \d_HADDR_0_iv_0_2[21]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_21_S, B => 
        \d_HADDR_0_iv_0_0[21]_net_1\, C => N_4514, D => N_247, Y
         => \d_HADDR_0_iv_0_2[21]_net_1\);
    
    \d_acc_1_0[7]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_789, B => \d_acc_1_0_0[7]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(7), Y => \d_acc[7]\);
    
    \state_RNICLIN[22]\ : CFG3
      generic map(INIT => x"23")

      port map(A => \state[22]_net_1\, B => N_290, C => N_272, Y
         => N_542_2);
    
    \d_acc_1[0]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_789, B => \d_acc_1_0[0]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(0), Y => \d_acc[0]\);
    
    \state[8]\ : SLE
      port map(D => \state_ns[20]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[8]_net_1\);
    
    un13_d_haddr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[8]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_5\, S => un13_d_haddr_1_cry_6_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_6\);
    
    \d_acc_1_0[18]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[18]_net_1\, B => \acc[18]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[18]_net_1\);
    
    un1_state_44_0_a3_2 : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \state[0]_net_1\, B => \pause_count[4]_net_1\, 
        C => \pause_count[3]_net_1\, D => N_4811, Y => N_4855);
    
    \haddr_fetch[11]\ : SLE
      port map(D => N_119_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[11]_net_1\);
    
    \haddr_write[23]\ : SLE
      port map(D => un46_d_haddr_cry_23_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[23]_net_1\);
    
    \envm_soft_reset[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_696_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \envm_soft_reset[0]_net_1\);
    
    \mask[13]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(13), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[13]_net_1\);
    
    \HWDATA_int_RNO_0[28]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_278, C => 
        \acc[28]_net_1\, D => \rdata[12]_net_1\, Y => 
        d_HWDATA_0_iv_2_1532_5_0);
    
    \d_ins2[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(9), B => un28_opcode, 
        Y => \d_ins2[9]_net_1\);
    
    \mask[18]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(18), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[18]_net_1\);
    
    \d_acc_1_0[3]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[3]_net_1\, B => \acc[3]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[3]_net_1\);
    
    \rdata[20]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(20), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[20]_net_1\);
    
    \HADDR_int[0]\ : SLE
      port map(D => \d_HADDR[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[0]\);
    
    \d_HADDR_0_iv_0[21]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[21]_net_1\, C => 
        \haddr_fetch[21]_net_1\, Y => \d_HADDR[21]\);
    
    \count_RNO_2[1]\ : CFG4
      generic map(INIT => x"0233")

      port map(A => N_252, B => d_N_3_mux_0, C => N_294, D => 
        \d_count_0_o2_0_1_2[1]\, Y => N_445);
    
    \ins1[17]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(17), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[17]_net_1\);
    
    \HWDATA_int[29]\ : SLE
      port map(D => \HWDATA_int_RNO[29]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(29));
    
    \state[22]\ : SLE
      port map(D => N_170, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[22]_net_1\);
    
    \d_HADDR_0_iv_1_0[1]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_1[1]_net_1\, B => 
        \haddr_fetch[1]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1_0[1]_net_1\);
    
    \HADDR_int[27]\ : SLE
      port map(D => \d_HADDR[27]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[27]\);
    
    \acc[22]\ : SLE
      port map(D => \d_acc[22]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[22]_net_1\);
    
    \haddr_fetch_RNO[2]\ : CFG3
      generic map(INIT => x"56")

      port map(A => \ConfigMaster_0_M_HADDR[2]\, B => N_4812, C
         => N_198, Y => N_64_i);
    
    \count_RNO_7[1]\ : CFG4
      generic map(INIT => x"F0F2")

      port map(A => \count[1]_net_1\, B => \state[22]_net_1\, C
         => \d_count_0_a2_2_0[1]\, D => N_259, Y => 
        \d_count_0_0_tz[1]\);
    
    state_m3_i_4 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[2]_net_1\, B => \state[5]_net_1\, C
         => \state_ns[22]\, D => \state_m3_i_2\, Y => 
        \state_m3_i_4\);
    
    \HWDATA_int_RNO_2[15]\ : CFG4
      generic map(INIT => x"FFF2")

      port map(A => N_2573_1, B => N_252, C => 
        d_HWDATA_0_iv_15_992_0, D => N_2063, Y => 
        d_HWDATA_0_iv_15_992_2);
    
    \d_HADDR_0_iv_2_RNO[20]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[20]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[20]\);
    
    \haddr_fetch[10]\ : SLE
      port map(D => N_4364_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[10]_net_1\);
    
    \expected[13]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(13), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[13]_net_1\);
    
    \count_RNO_4[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_541, B => N_266, C => 
        \d_count_0_a2_1_2_1[1]\, Y => \d_count_0_a2_1_c_1[1]\);
    
    un7_hready_2_RNI8KKE : CFG4
      generic map(INIT => x"0800")

      port map(A => \count[1]_net_1\, B => un9_hready_2, C => 
        \ins1[21]_net_1\, D => \ins1[20]_net_1\, Y => N_591);
    
    d_count_1_sqmuxa_i_a2_0_o2_i_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \state[23]_net_1\, B => \state[24]_net_1\, Y
         => N_259);
    
    \HWDATA_int_RNO[0]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => d_HWDATA_0_iv_30_380_1_0, B => N_178, C => 
        d_HWDATA_0_iv_30_380_1_2, Y => \HWDATA_int_RNO[0]_net_1\);
    
    \state[1]\ : SLE
      port map(D => \state[2]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[1]_net_1\);
    
    \haddr_write[4]\ : SLE
      port map(D => un46_d_haddr_cry_4_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[4]_net_1\);
    
    \HADDR_int[28]\ : SLE
      port map(D => \d_HADDR[28]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[28]\);
    
    \bytecount[7]\ : SLE
      port map(D => N_40_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[7]_net_1\);
    
    \d_HADDR_0_iv_0_a2_3[0]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[0]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4764);
    
    un22_opcode_0_0_a2 : CFG4
      generic map(INIT => x"001A")

      port map(A => \ins1[26]_net_1\, B => \ins1[24]_net_1\, C
         => \ins1[25]_net_1\, D => N_80, Y => N_97);
    
    \mask[26]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(26), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[26]_net_1\);
    
    \d_HADDR_0_iv_0[4]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => un13_d_haddr_1_cry_2_S, B => \state[5]_net_1\, 
        C => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0[4]_net_1\);
    
    \acc[13]\ : SLE
      port map(D => \d_acc[13]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[13]_net_1\);
    
    \HWDATA_int[7]\ : SLE
      port map(D => \HWDATA_int_RNO[7]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(7));
    
    \rdata[7]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(7), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[7]_net_1\);
    
    \bytecount_RNO[7]\ : CFG3
      generic map(INIT => x"70")

      port map(A => \state[21]_net_1\, B => N_109_i, C => N_108, 
        Y => N_40_i_0);
    
    \ins1[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[0]_net_1\);
    
    un46_d_haddr_cry_0_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \HADDR_int_fast[0]_net_1\, B => 
        \ins1[16]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        GND_net_1, S => OPEN, Y => OPEN, FCO => 
        un46_d_haddr_cry_0_0_FCO);
    
    \d_HADDR_0_iv_1[14]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_0[14]_net_1\, B => 
        \haddr_fetch[14]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1[14]_net_1\);
    
    \rdata_RNIE9J21[21]\ : CFG4
      generic map(INIT => x"33B3")

      port map(A => \state[21]_net_1\, B => N_4885, C => 
        \rdata[21]_net_1\, D => \count[0]_net_1\, Y => 
        d_HWDATA_0_iv_25_605_7_1_0);
    
    \HWDATA_int[17]\ : SLE
      port map(D => \HWDATA_int_RNO[17]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(17));
    
    un7_hready_2 : CFG2
      generic map(INIT => x"1")

      port map(A => \ins1[22]_net_1\, B => \ins1[23]_net_1\, Y
         => un9_hready_2);
    
    \HADDR_int[19]\ : SLE
      port map(D => \d_HADDR[19]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[19]\);
    
    un1_state_25_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \state[7]_net_1\, B => \state[8]_net_1\, Y
         => N_789);
    
    \state_RNIUR1F[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => \state[26]_net_1\, Y => 
        N_700_i_0);
    
    \d_ins2[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(11), B => un28_opcode, 
        Y => \d_ins2[11]_net_1\);
    
    \state[24]\ : SLE
      port map(D => N_12_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[24]_net_1\);
    
    \HWDATA_int_RNO_3[25]\ : CFG4
      generic map(INIT => x"B3A0")

      port map(A => \state[10]_net_1\, B => N_263, C => 
        \acc[25]_net_1\, D => \rdata[9]_net_1\, Y => 
        d_HWDATA_0_iv_5_1424_0);
    
    \d_HADDR_0_iv_1[27]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[27]_net_1\, B => 
        \ins2[27]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_1[27]_net_1\);
    
    \d_HADDR_0_iv[31]\ : CFG4
      generic map(INIT => x"FCF8")

      port map(A => \un1_state_30_0_0\, B => 
        un13_d_haddr_1_s_29_S, C => \d_HADDR_0_iv_1_1[31]_net_1\, 
        D => N_4814, Y => \d_HADDR[31]\);
    
    \HADDR_int_RNO_0[3]\ : CFG4
      generic map(INIT => x"4445")

      port map(A => \d_HADDR_0_iv_0_0[3]_net_1\, B => 
        \haddr_fetch[3]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => \d_HADDR_0_iv_i_1[3]\);
    
    un7_hready_2_RNI7JKE : CFG4
      generic map(INIT => x"AE2A")

      port map(A => \count[0]_net_1\, B => un9_hready_2, C => 
        \ins1[21]_net_1\, D => \ins1[20]_net_1\, Y => N_276);
    
    \haddr_fetch[6]\ : SLE
      port map(D => N_4720_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[6]_net_1\);
    
    \bytecount_RNIDL3T[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \bytecount[0]_net_1\, B => 
        \bytecount[1]_net_1\, Y => N_266);
    
    \haddr_fetch[27]\ : SLE
      port map(D => N_4407_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[27]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_2_0_0 : CFG4
      generic map(INIT => x"A8EC")

      port map(A => \state[16]_net_1\, B => N_117, C => 
        d_state61_li, D => HREADY_i_3, Y => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\);
    
    un1_rdata_0_I_80_i_x2_0 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[16]_net_1\, B => \rdata[16]_net_1\, 
        C => \mask[16]_net_1\, Y => N_323_i);
    
    un1_rdata_0_I_69 : ARI1
      generic map(INIT => x"40095")

      port map(A => un1_rdata_0_N_22, B => \expected[30]_net_1\, 
        C => \mask[30]_net_1\, D => \rdata[30]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[14]\, S => OPEN, Y => OPEN, FCO => 
        d_state61_li);
    
    \HWDATA_int_RNO_0[26]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_4_1460_5_0, B => N_4577, C => 
        \rdata[26]_net_1\, D => N_403, Y => 
        d_HWDATA_0_iv_4_1460_5_2);
    
    pause_count_n2_i_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \pause_count[2]_net_1\, B => 
        \pause_count[1]_net_1\, C => \pause_count[0]_net_1\, Y
         => N_66_i);
    
    \HADDR_int[20]\ : SLE
      port map(D => \d_HADDR[20]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[20]\);
    
    un1_d_HWRITE_0_sqmuxa_5_i_a2 : CFG3
      generic map(INIT => x"08")

      port map(A => \state[21]_net_1\, B => N_109_i, C => 
        HREADY_i_3, Y => N_212);
    
    \haddr_write[14]\ : SLE
      port map(D => un46_d_haddr_cry_14_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[14]_net_1\);
    
    \HWDATA_int_RNO_1[22]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \rdata[6]_net_1\, B => \count[1]_net_1\, C
         => N_274, D => N_252, Y => N_4653);
    
    \haddr_fetch_RNO[7]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_5_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[7]\, D => N_4812, Y => 
        \haddr_fetch_RNO[7]_net_1\);
    
    \d_acc_1_0[28]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[28]_net_1\, B => \acc[28]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[28]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa : CFG4
      generic map(INIT => x"FCEC")

      port map(A => \d_HWRITE_0_sqmuxa_1_0_a3_1\, B => 
        d_HWRITE_0_sqmuxa_2, C => \un1_d_HWRITE_0_sqmuxa_0_2\, D
         => \d_HTRANS_0_sqmuxa_4_1\, Y => \un1_d_HWRITE_0_sqmuxa\);
    
    \d_HADDR_0_iv_0_0[16]\ : CFG4
      generic map(INIT => x"5703")

      port map(A => un13_d_haddr_1_cry_14_S, B => 
        \haddr_write[16]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[16]_net_1\);
    
    \pause_count_RNO[1]\ : CFG4
      generic map(INIT => x"006F")

      port map(A => \pause_count[0]_net_1\, B => 
        \pause_count[1]_net_1\, C => N_4813, D => N_3400, Y => 
        N_37_i_0);
    
    \pause_count[0]\ : SLE
      port map(D => N_4316_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        pause_counte, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pause_count[0]_net_1\);
    
    un46_d_haddr_cry_27 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[27]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_26\, S => un46_d_haddr_cry_27_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_27\);
    
    un46_d_haddr_cry_23 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[23]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_22\, S => un46_d_haddr_cry_23_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_23\);
    
    \state_ns_0[8]\ : CFG4
      generic map(INIT => x"FAFE")

      port map(A => \state_ns_0_0[8]_net_1\, B => 
        \state_ns_0_a3_2[8]_net_1\, C => N_186, D => HREADY_i_3, 
        Y => \state_ns[8]\);
    
    un13_d_haddr_1_cry_23 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[25]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_22\, S => un13_d_haddr_1_cry_23_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_23\);
    
    d_HWRITE_0_sqmuxa_4_0 : CFG3
      generic map(INIT => x"FE")

      port map(A => N_404, B => N_402, C => N_403, Y => 
        d_HWRITE_0_sqmuxa_4);
    
    \mask[27]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(27), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[27]_net_1\);
    
    \haddr_write[1]\ : SLE
      port map(D => un46_d_haddr_cry_1_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[1]_net_1\);
    
    \HWDATA_int[14]\ : SLE
      port map(D => \HWDATA_int_RNO[14]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(14));
    
    \bytecount_RNO[11]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4340, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_48_i_0);
    
    state_21_rep1_RNI7JG7O : CFG4
      generic map(INIT => x"EECE")

      port map(A => \state_21_rep1\, B => 
        un1_state_31_i_i_a2_0_d_0_0_0, C => 
        \un1_state_31_i_i_a2_0_d_0_0_1\, D => 
        un1_state_31_i_i_a2_0_d_1_0_1, Y => N_164);
    
    un46_d_haddr_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[7]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_6\, S => un46_d_haddr_cry_7_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_7\);
    
    \d_HADDR_0_iv_0_0[13]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => un13_d_haddr_1_cry_11_S, B => \state_ns[0]\, 
        C => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0_0[13]_net_1\);
    
    \rdata_RNI00L91[16]\ : CFG4
      generic map(INIT => x"F2FF")

      port map(A => \count[1]_net_1\, B => \rdata[16]_net_1\, C
         => N_465, D => N_251, Y => 
        d_HWDATA_0_iv_14_1028_2_a2_i_1);
    
    \HADDR_int_RNO[3]\ : CFG4
      generic map(INIT => x"5040")

      port map(A => \d_HADDR_0_iv_0_2[3]_net_1\, B => 
        un46_d_haddr_cry_3_S, C => \d_HADDR_0_iv_i_1[3]\, D => 
        N_247, Y => \d_HADDR_0_iv_i_0[3]\);
    
    un46_d_haddr_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[4]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_3\, S => un46_d_haddr_cry_4_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_4\);
    
    d_HADDR_0_sqmuxa_1_i_a2_0_a3_0_a2_RNIJMHRN : CFG4
      generic map(INIT => x"FFFE")

      port map(A => defSlaveSMNextState_m_0_2, B => N_837, C => 
        un1_state_31_i_i_a2_0_d_1_0_1, D => 
        defSlaveSMNextState_m_0_3, Y => N_4873);
    
    un46_d_haddr_cry_28 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[28]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_27\, S => un46_d_haddr_cry_28_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_28\);
    
    \acc[18]\ : SLE
      port map(D => \d_acc[18]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[18]_net_1\);
    
    un13_d_haddr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[6]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_3\, S => un13_d_haddr_1_cry_4_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_4\);
    
    d_HADDR_0_sqmuxa_1_i_a2_0_a3_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \state[24]_net_1\, B => \state[14]_net_1\, C
         => \state[19]_net_1\, D => \state[11]_net_1\, Y => N_837);
    
    d_count_1_sqmuxa_i_a2_0_o2_i_o2_RNIS4TE : CFG2
      generic map(INIT => x"D")

      port map(A => N_272, B => N_259, Y => N_369);
    
    \count_RNI2UJ11[0]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => \state[21]_net_1\, B => N_403, C => 
        \count[0]_net_1\, Y => d_HWDATA_0_iv_7_1343_o2_0_0);
    
    \d_acc_1[13]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[13]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(13), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[13]\);
    
    un1_state_39_2_i_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[10]_net_1\, B => \state[4]_net_1\, Y
         => N_200);
    
    \haddr_fetch[12]\ : SLE
      port map(D => N_4402_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[12]_net_1\);
    
    \HADDR_int[1]\ : SLE
      port map(D => \d_HADDR[1]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[1]\);
    
    un46_d_haddr_cry_30_3 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[11]\, B => 
        \ConfigMaster_0_M_HADDR[8]\, C => 
        \ConfigMaster_0_M_HADDR[9]\, D => 
        \ConfigMaster_0_M_HADDR[10]\, FCI => 
        un46_d_haddr_cry_30_1_FCO, S => OPEN, Y => OPEN, FCO => 
        un46_d_haddr_cry_30_3_FCO);
    
    \d_HADDR_0_iv_0_a2_3[16]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \ins2[16]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4759);
    
    \haddr_write[11]\ : SLE
      port map(D => un46_d_haddr_cry_11_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[11]_net_1\);
    
    \d_HADDR_0_iv_0_a2_0[7]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => un13_d_haddr_1_cry_5_S, B => 
        \un1_state_30_0_0\, C => N_4814, Y => N_4592);
    
    \rdata_RNIOIFC1[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_600, B => \rdata[9]_net_1\, Y => N_582);
    
    un46_d_haddr_cry_1_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[17]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[1]\, C => GND_net_1, D => 
        GND_net_1, FCI => un46_d_haddr_cry_0_0_FCO, S => OPEN, Y
         => OPEN, FCO => un46_d_haddr_cry_1_0_FCO);
    
    \state_ns_i_a2_10_i_1[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \ins1[31]_net_1\, B => \state[4]_net_1\, C
         => \state[3]_net_1\, Y => 
        \state_ns_i_a2_10_i_1[1]_net_1\);
    
    \d_acc[9]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1146, C => 
        \ins2[9]_net_1\, D => \acc[9]_net_1\, Y => 
        \d_acc[9]_net_1\);
    
    un13_d_haddr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[11]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_8\, S => un13_d_haddr_1_cry_9_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_9\);
    
    \acc[31]\ : SLE
      port map(D => \d_acc[31]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[31]_net_1\);
    
    \rdata[17]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(17), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[17]_net_1\);
    
    \HADDR_int_RNO[30]\ : CFG4
      generic map(INIT => x"5040")

      port map(A => \d_HADDR_0_iv_0_2[30]_net_1\, B => 
        un46_d_haddr_cry_30_S, C => \d_HADDR_0_iv_i_1[30]\, D => 
        N_247, Y => \d_HADDR_0_iv_i_0[30]\);
    
    \expected[23]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(23), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[23]_net_1\);
    
    \d_HADDR_0_iv_0_0[17]\ : CFG4
      generic map(INIT => x"5703")

      port map(A => un13_d_haddr_1_cry_15_S, B => 
        \haddr_write[17]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[17]_net_1\);
    
    \ins2[1]\ : SLE
      port map(D => \d_ins2[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[1]_net_1\);
    
    \haddr_fetch_RNO[28]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_26_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[28]\, D => N_4812, Y => N_19_i_0);
    
    \d_HADDR_0_iv_RNO[29]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => un13_d_haddr_1_cry_27_S, B => 
        \un1_state_30_0_0\, C => N_4814, Y => 
        \un13_d_haddr_1_m[29]\);
    
    \ins2[7]\ : SLE
      port map(D => \d_ins2[7]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[7]_net_1\);
    
    \HWDATA_int_RNO_0[5]\ : CFG4
      generic map(INIT => x"CCEC")

      port map(A => N_252, B => d_HWDATA_0_iv_25_605_7_0, C => 
        N_4541, D => N_274, Y => d_HWDATA_0_iv_25_605_7_1);
    
    \state_RNIVR0F[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => \state[18]_net_1\, Y => 
        N_702_i_0);
    
    \d_HADDR_0_iv_1[29]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[29]_net_1\, B => 
        \ins2[29]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_1[29]_net_1\);
    
    \count_RNIGI2A[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \count[1]_net_1\, B => \state[21]_net_1\, Y
         => N_263);
    
    \count_RNI1TLE[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_4916, B => \count[1]_net_1\, Y => N_592);
    
    \ins1[3]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(3), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[3]_net_1\);
    
    \HWDATA_int_RNO_0[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[10]_net_1\, D => \rdata[26]_net_1\, Y => 
        d_HWDATA_0_iv_20_812_0_0);
    
    \rdata[5]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(5), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[5]_net_1\);
    
    \bytecount[2]\ : SLE
      port map(D => N_32_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[2]_net_1\);
    
    \HWDATA_int_RNO_2[31]\ : CFG3
      generic map(INIT => x"13")

      port map(A => \state[10]_net_1\, B => N_2066, C => 
        \acc[31]_net_1\, Y => d_HWDATA_0_iv_1640_2_1);
    
    \d_acc_1_0[10]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[10]_net_1\, B => \acc[10]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[10]_net_1\);
    
    \HWDATA_int_RNO_0[15]\ : CFG3
      generic map(INIT => x"80")

      port map(A => d_HWDATA_0_iv_1640_a8_3_0, B => N_276, C => 
        \count[1]_net_1\, Y => N_2060);
    
    \count_RNO_0[1]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => d_m2_e_2_2, B => N_375, C => 
        \d_count_0_a2_1_2_1[1]\, D => N_541, Y => 
        \d_count_0_a2_1_d[1]\);
    
    \rdata_RNIPV3M[24]\ : CFG4
      generic map(INIT => x"53FF")

      port map(A => \rdata[24]_net_1\, B => \rdata[8]_net_1\, C
         => \count[1]_net_1\, D => N_249, Y => 
        d_HWDATA_0_iv_14_1028_0_a2_i_1);
    
    un46_d_haddr_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[19]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[3]\, C => GND_net_1, D => 
        GND_net_1, FCI => \un46_d_haddr_cry_2\, S => 
        un46_d_haddr_cry_3_S, Y => OPEN, FCO => 
        \un46_d_haddr_cry_3\);
    
    un13_d_haddr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[5]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_2\, S => un13_d_haddr_1_cry_3_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_3\);
    
    \state_ns_i_a2_10_i_2[1]\ : CFG4
      generic map(INIT => x"AABA")

      port map(A => \state_ns_i_a2_10_i_1[1]_net_1\, B => 
        \state[9]_net_1\, C => N_138, D => N_789, Y => 
        \state_ns_i_a2_10_i_2[1]_net_1\);
    
    \ins1[19]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(19), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[19]_net_1\);
    
    busy : SLE
      port map(D => d_busy, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \state[2]_net_1\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \busy\);
    
    \d_HADDR_0_iv_1_0[22]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_1[22]_net_1\, B => 
        \haddr_fetch[22]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1_0[22]_net_1\);
    
    un4_bytecount_0_o2_i_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => d_N_3_mux_0, B => N_266, Y => N_109_i);
    
    \d_acc_0[6]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[6]_net_1\, B => \ins2[6]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(6), D => \state[8]_net_1\, Y => 
        N_1143);
    
    \expected[8]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(8), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[8]_net_1\);
    
    \un7_iv[14]\ : CFG4
      generic map(INIT => x"F0FD")

      port map(A => \un7_iv_1[14]_net_1\, B => 
        un1_state_31_i_i_a2_0_d_1_0_1, C => un1_state_31_i_i_o2_0, 
        D => \un7_iv_0_a1_0[14]_net_1\, Y => \un7_iv[14]_net_1\);
    
    \HWDATA_int[16]\ : SLE
      port map(D => \HWDATA_int_RNO[16]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(16));
    
    \bytecount[14]\ : SLE
      port map(D => N_55_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[14]_net_1\);
    
    \d_ins2[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(21), B => un28_opcode, 
        Y => \d_ins2[21]_net_1\);
    
    \rdata[31]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(31), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[31]_net_1\);
    
    \d_ins2[19]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(19), B => un28_opcode, 
        Y => \d_ins2[19]_net_1\);
    
    \acc[15]\ : SLE
      port map(D => \d_acc[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[15]_net_1\);
    
    \state_ns_0_a3_2_3[8]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \state[16]_net_1\, B => \state[15]_net_1\, C
         => \ins1[31]_net_1\, D => \state[14]_net_1\, Y => 
        \state_ns_0_a3_2_3[8]_net_1\);
    
    un1_state_46_3 : CFG4
      generic map(INIT => x"FDEC")

      port map(A => HREADY_i_3, B => \un1_state_46_1\, C => N_789, 
        D => \un1_state_39\, Y => \un1_state_46_3\);
    
    \bytecount[11]\ : SLE
      port map(D => N_48_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[11]_net_1\);
    
    \haddr_write[16]\ : SLE
      port map(D => un46_d_haddr_cry_16_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[16]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_0_2 : CFG3
      generic map(INIT => x"80")

      port map(A => \un12_size_2_0_5\, B => \un12_size_2_0_4\, C
         => \un1_d_HWRITE_0_sqmuxa_0_1\, Y => 
        \un1_d_HWRITE_0_sqmuxa_0_2\);
    
    \d_HADDR_0_iv_1[4]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_0[4]_net_1\, B => 
        \haddr_fetch[4]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1[4]_net_1\);
    
    \count_RNIOP5V2[1]\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \d_count_0_o2_0[1]\, B => HREADY_i_3, C => 
        \count[1]_net_1\, D => N_281, Y => N_319);
    
    \state_RNO[27]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_148, B => \state_m3_i_8\, C => N_101, D => 
        \state_m3_i_a3\, Y => N_741_i_0);
    
    \haddr_fetch[8]\ : SLE
      port map(D => N_4365_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[8]_net_1\);
    
    \d_ins2[30]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(30), B => un28_opcode, 
        Y => \d_ins2[30]_net_1\);
    
    \state_ns_0_o2[7]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \state[22]_net_1\, B => \state[21]_net_1\, C
         => HREADY_i_3, Y => N_101);
    
    d_HWDATA_0_sqmuxa_2 : CFG4
      generic map(INIT => x"AAA8")

      port map(A => \state[21]_net_1\, B => N_109_i, C => 
        defSlaveSMNextState_m, D => \un1_hready_2_0_0\, Y => 
        \d_HWDATA_0_sqmuxa_2\);
    
    \acc[16]\ : SLE
      port map(D => \d_acc[16]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[16]_net_1\);
    
    \HWDATA_int[11]\ : SLE
      port map(D => N_1926, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(11));
    
    \state_ns_i_a2_13_0_a3_5[1]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \state[26]_net_1\, B => \state[20]_net_1\, C
         => \state_ns_i_a2_13_0_a3_5_0[1]_net_1\, D => 
        \un1_state_39_3\, Y => \state_ns_i_a2_13_0_a3_5[1]_net_1\);
    
    \state_ns_0[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \state_ns_0_a2_0_1[5]_net_1\, B => HREADY_i_3, 
        C => \state[23]_net_1\, Y => \state_ns[5]\);
    
    \bytecount_RNI6N7Q1[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \bytecount[5]_net_1\, B => 
        \bytecount[4]_net_1\, C => \bytecount[3]_net_1\, D => 
        \bytecount[2]_net_1\, Y => d_m1_e_1_1);
    
    \d_HADDR_0_iv_0[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[0]_net_1\, C => \haddr_fetch[0]_net_1\, 
        Y => \d_HADDR[0]\);
    
    \d_acc_0[11]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[11]_net_1\, B => \ins2[11]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(11), D => \state[8]_net_1\, Y => 
        N_1148);
    
    \state_RNIHJ2A[22]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \count[1]_net_1\, B => \state[22]_net_1\, Y
         => N_4711);
    
    \state_fast[21]\ : SLE
      port map(D => \state_ns_fast[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \state_fast[21]_net_1\);
    
    \haddr_fetch[1]\ : SLE
      port map(D => \ConfigMaster_0_M_HADDR[1]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[1]_net_1\);
    
    un13_d_haddr_1_cry_25 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[27]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_24\, S => un13_d_haddr_1_cry_25_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_25\);
    
    \state_ns_i_o2_0[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_4855, B => N_3400, Y => \state_ns[28]\);
    
    un13_d_haddr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[15]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un13_d_haddr_1_cry_27_5_FCO, S => un13_d_haddr_1_cry_13_S, 
        Y => OPEN, FCO => \un13_d_haddr_1_cry_13\);
    
    \state_RNIHJ2A_0[22]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \count[1]_net_1\, B => \state[22]_net_1\, Y
         => \d_count_0_a3_8_0[1]\);
    
    un1_rdata_0_I_92_i_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[2]_net_1\, B => \rdata[2]_net_1\, C
         => \mask[2]_net_1\, Y => N_347_i);
    
    \state[0]\ : SLE
      port map(D => \state_ns[28]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[0]_net_1\);
    
    un46_d_haddr_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[17]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[1]\, C => GND_net_1, D => 
        GND_net_1, FCI => \un46_d_haddr_cry_0\, S => 
        un46_d_haddr_cry_1_S, Y => OPEN, FCO => 
        \un46_d_haddr_cry_1\);
    
    \rdata[29]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(29), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[29]_net_1\);
    
    \d_HADDR_0_iv_0[6]\ : CFG4
      generic map(INIT => x"DDDC")

      port map(A => un13_d_haddr_1_cry_4_S, B => \state_ns[0]\, C
         => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0[6]_net_1\);
    
    \d_acc_1_0_0[7]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[7]_net_1\, B => \acc[7]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0_0[7]_net_1\);
    
    \d_acc[1]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1138, C => 
        \ins2[1]_net_1\, D => \acc[1]_net_1\, Y => 
        \d_acc[1]_net_1\);
    
    \rdata[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[0]_net_1\);
    
    \HADDR_int[17]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[17]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[17]\);
    
    \HWDATA_int_RNO_0[0]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => \state[10]_net_1\, B => N_4889, C => 
        \acc[0]_net_1\, Y => d_HWDATA_0_iv_30_380_1_0);
    
    un1_d_HWRITE_1_sqmuxa_2_i_a2_0_0 : CFG3
      generic map(INIT => x"80")

      port map(A => N_249, B => d_N_3_mux_0, C => 
        \d_HWRITE_1_sqmuxa_1_i_a2_0_a2_0\, Y => 
        \un1_d_HWRITE_1_sqmuxa_2_i_a2_0_0\);
    
    \count_RNO_8[0]\ : CFG4
      generic map(INIT => x"A022")

      port map(A => \count[0]_net_1\, B => N_259, C => N_290, D
         => N_251, Y => N_543);
    
    un46_d_haddr_cry_22 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[22]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_21\, S => un46_d_haddr_cry_22_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_22\);
    
    \count[0]\ : SLE
      port map(D => N_4888_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \count[0]_net_1\);
    
    \rdata_RNIK9US1[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[18]_net_1\, B => \rdata[2]_net_1\, C
         => N_592, D => N_254, Y => N_4556_1);
    
    \HWDATA_int[10]\ : SLE
      port map(D => N_1897, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(10));
    
    \d_acc_0[27]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[27]_net_1\, B => \ins2[27]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(27), D => \state[8]_net_1\, Y => 
        N_1164);
    
    \d_acc[17]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1154, C => 
        \ins2[17]_net_1\, D => \acc[17]_net_1\, Y => 
        \d_acc[17]_net_1\);
    
    \state[21]\ : SLE
      port map(D => \state_ns[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[21]_net_1\);
    
    \ins1_RNIUCDVT3[5]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[5]_net_1\, B => N_78, C => N_164, 
        D => \ins1[5]_net_1\, FCI => d_bytecount_i_m2_cry_4, S
         => N_106, Y => OPEN, FCO => d_bytecount_i_m2_cry_5);
    
    un13_d_haddr_1_cry_28 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[30]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_27\, S => un13_d_haddr_1_cry_28_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_28\);
    
    \mask[31]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(31), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[31]_net_1\);
    
    \rdata_RNIJ9VS1[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[22]_net_1\, B => \rdata[6]_net_1\, C
         => N_592, D => N_254, Y => N_680_2);
    
    \haddr_fetch[25]\ : SLE
      port map(D => N_3162_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[25]_net_1\);
    
    \count_RNI91JR[0]\ : CFG4
      generic map(INIT => x"7F3F")

      port map(A => \count[0]_net_1\, B => N_251, C => N_252, D
         => N_249, Y => N_291);
    
    \bytecount_RNO[10]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4339, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_46_i_0);
    
    \acc[5]\ : SLE
      port map(D => \d_acc[5]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[5]_net_1\);
    
    \acc[11]\ : SLE
      port map(D => \d_acc[11]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[11]_net_1\);
    
    un46_d_haddr_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[8]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_7\, S => un46_d_haddr_cry_8_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_8\);
    
    un1_state_30_0 : CFG2
      generic map(INIT => x"E")

      port map(A => N_4814, B => \un1_state_30_0_0\, Y => 
        un1_state_30);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => defSlaveSMNextState_m_0_2, B => 
        \un1_d_HWRITE_1_sqmuxa_2_i_o3_0\, C => 
        un1_state_31_i_i_a2_0_d_1_0_1, D => 
        defSlaveSMNextState_m_0_3, Y => N_294);
    
    \haddr_write[28]\ : SLE
      port map(D => un46_d_haddr_cry_28_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[28]_net_1\);
    
    \haddr_fetch_RNO[25]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_23_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[25]\, D => N_4812, Y => 
        N_3162_i_0);
    
    \d_HADDR_0_iv_0[13]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_0_2[13]_net_1\, B => 
        un46_d_haddr_cry_13_S, C => \d_HADDR_0_iv_0_1[13]_net_1\, 
        D => N_247, Y => \d_HADDR[13]\);
    
    \state_RNIS2GD[22]\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_252, B => \state[22]_net_1\, Y => N_317);
    
    \bytecount[0]\ : SLE
      port map(D => N_28_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[0]_net_1\);
    
    \d_HADDR_0_iv_0_2[18]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_18_S, B => 
        \d_HADDR_0_iv_0_0[18]_net_1\, C => N_4387, D => N_247, Y
         => \d_HADDR_0_iv_0_2[18]_net_1\);
    
    \state[12]\ : SLE
      port map(D => \state_ns[16]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[12]_net_1\);
    
    \state_RNIBKIN_0[22]\ : CFG4
      generic map(INIT => x"C8C0")

      port map(A => \state[22]_net_1\, B => \count[0]_net_1\, C
         => \state[21]_net_1\, D => N_252, Y => 
        d_HWDATA_0_iv_20_812_o3_0_0);
    
    \ins1[10]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(10), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[10]_net_1\);
    
    \HADDR_int[18]\ : SLE
      port map(D => \d_HADDR[18]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[18]\);
    
    \mask[24]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(24), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[24]_net_1\);
    
    \mask[15]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(15), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[15]_net_1\);
    
    \bytecount[10]\ : SLE
      port map(D => N_46_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[10]_net_1\);
    
    \state_RNIRAVI[22]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \state[21]_net_1\, B => \state[22]_net_1\, Y
         => N_251);
    
    \ins2[3]\ : SLE
      port map(D => \d_ins2[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[3]_net_1\);
    
    \count_RNIFK6P1[1]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \count[1]_net_1\, B => N_403, C => N_258, Y
         => N_270);
    
    \d_HADDR_0_iv_0_0[24]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_0_0_0[24]_net_1\, B => 
        un46_d_haddr_cry_24_S, C => 
        \d_HADDR_0_iv_0_0_1[24]_net_1\, D => N_247, Y => 
        \d_HADDR[24]\);
    
    \d_bytecount_RNO[15]\ : ARI1
      generic map(INIT => x"4D782")

      port map(A => \ins1[15]_net_1\, B => N_78, C => N_164, D
         => \bytecount[15]_net_1\, FCI => d_bytecount_i_m2_cry_14, 
        S => N_1116, Y => OPEN, FCO => OPEN);
    
    un46_d_haddr_cry_16 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[16]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un46_d_haddr_cry_30_5_FCO, S => un46_d_haddr_cry_16_S, Y
         => OPEN, FCO => \un46_d_haddr_cry_16\);
    
    \d_acc_1[4]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[4]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(4), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[4]\);
    
    \rdata_RNIB5142[8]\ : CFG4
      generic map(INIT => x"FBF0")

      port map(A => N_263, B => \rdata[8]_net_1\, C => 
        d_HWDATA_0_iv_14_1028_2_a2_i_1, D => N_249, Y => N_4889);
    
    \HWDATA_int_RNO_0[19]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_601, C => 
        \acc[19]_net_1\, D => \rdata[3]_net_1\, Y => 
        d_HWDATA_0_iv_11_1163_0_0);
    
    \d_acc[19]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1156, C => 
        \ins2[19]_net_1\, D => \acc[19]_net_1\, Y => 
        \d_acc[19]_net_1\);
    
    \count_RNIJHMB1[0]\ : CFG4
      generic map(INIT => x"F2F3")

      port map(A => \state[21]_net_1\, B => \count[0]_net_1\, C
         => N_403, D => N_4711, Y => N_4625);
    
    \HWDATA_int_RNO[17]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \rdata[1]_net_1\, B => N_601, C => 
        d_HWDATA_0_iv_13_1073_0_1, D => N_296, Y => 
        \HWDATA_int_RNO[17]_net_1\);
    
    \HWDATA_int_RNO_4[25]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \count[1]_net_1\, B => \rdata[25]_net_1\, Y
         => d_HWDATA_0_iv_5_1424_a8_0_0);
    
    \d_acc_1[18]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[18]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(18), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[18]\);
    
    \HWDATA_int_RNO_0[20]\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => N_512_1, B => N_4625, C => \rdata[20]_net_1\, 
        D => N_485, Y => d_HWDATA_0_iv_10_1208_0_1);
    
    \haddr_write[19]\ : SLE
      port map(D => un46_d_haddr_cry_19_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[19]_net_1\);
    
    \d_acc[2]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1139, C => 
        \ins2[2]_net_1\, D => \acc[2]_net_1\, Y => 
        \d_acc[2]_net_1\);
    
    \d_ins2[14]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(14), B => un28_opcode, 
        Y => \d_ins2[14]_net_1\);
    
    \d_acc[23]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1160, C => 
        \ins2[23]_net_1\, D => \acc[23]_net_1\, Y => 
        \d_acc[23]_net_1\);
    
    \HWDATA_int_RNO_0[25]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \rdata[25]_net_1\, B => \state[22]_net_1\, C
         => N_252, D => d_HWDATA_0_iv_5_1424_0, Y => 
        d_HWDATA_0_iv_5_1424_1);
    
    \expected[17]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(17), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[17]_net_1\);
    
    \mask[30]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(30), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[30]_net_1\);
    
    un1_rdata_0_I_27 : ARI1
      generic map(INIT => x"40095")

      port map(A => un1_rdata_0_N_57, B => \expected[6]_net_1\, C
         => \mask[6]_net_1\, D => \rdata[6]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[2]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[3]\);
    
    \state_ns_0_0_a3[17]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => defSlaveSMNextState_m_0_2, B => 
        \state[25]_net_1\, C => un1_state_31_i_i_a2_0_d_1_0_1, D
         => defSlaveSMNextState_m_0_3, Y => N_654);
    
    \HWDATA_int_RNO[27]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \rdata[27]_net_1\, B => N_4777_1, C => 
        d_HWDATA_0_iv_3_1496_0_2, D => N_683_2, Y => 
        \HWDATA_int_RNO[27]_net_1\);
    
    pause_count_n3_i_o2 : CFG3
      generic map(INIT => x"7F")

      port map(A => \pause_count[2]_net_1\, B => 
        \pause_count[1]_net_1\, C => \pause_count[0]_net_1\, Y
         => N_4811);
    
    un13_d_haddr_1_cry_27_1 : ARI1
      generic map(INIT => x"48000")

      port map(A => \ConfigMaster_0_M_HADDR[6]\, B => 
        \ConfigMaster_0_M_HADDR[3]\, C => 
        \ConfigMaster_0_M_HADDR[4]\, D => 
        \ConfigMaster_0_M_HADDR[5]\, FCI => 
        \ConfigMaster_0_M_HADDR[2]\, S => OPEN, Y => OPEN, FCO
         => un13_d_haddr_1_cry_27_1_FCO);
    
    \ins1_RNIUC04_0[22]\ : CFG4
      generic map(INIT => x"FEFF")

      port map(A => \ins1[23]_net_1\, B => \ins1[22]_net_1\, C
         => \ins1[21]_net_1\, D => \ins1[20]_net_1\, Y => N_249);
    
    \haddr_fetch_RNO[5]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_3_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[5]\, D => N_4812, Y => 
        \haddr_fetch_RNO[5]_net_1\);
    
    \haddr_fetch[3]\ : SLE
      port map(D => N_53_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[3]_net_1\);
    
    d_HTRANS_0_sqmuxa_4_1 : CFG3
      generic map(INIT => x"02")

      port map(A => \bytecount[2]_net_1\, B => N_266, C => N_252, 
        Y => \d_HTRANS_0_sqmuxa_4_1\);
    
    \d_HADDR_0_iv_1_0[31]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => \d_HADDR_0_iv_1[31]_net_1\, B => 
        \haddr_fetch[31]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_1_0[31]_net_1\);
    
    \rdata_RNIFB9C2[21]\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => N_249, B => N_251, C => 
        d_HWDATA_0_iv_25_605_7_1_0, D => N_4472, Y => 
        d_HWDATA_0_iv_25_605_7_1_1);
    
    \d_acc_1_0[21]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[21]_net_1\, B => \acc[21]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[21]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_5_i_0_2 : CFG4
      generic map(INIT => x"0C08")

      port map(A => \un1_d_HWRITE_0_sqmuxa_5_i_a3_1_0\, B => 
        \state[21]_net_1\, C => HREADY_i_3, D => N_109_i, Y => 
        \un1_d_HWRITE_0_sqmuxa_5_i_0_2\);
    
    \HADDR_int[10]\ : SLE
      port map(D => \d_HADDR[10]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[10]\);
    
    un1_state_42_0_0_1 : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \state[28]_net_1\, B => \state[16]_net_1\, C
         => \state[6]_net_1\, D => N_125, Y => 
        \un1_state_42_0_0_1\);
    
    \count_RNO_2[0]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => \d_count_i_a2_1_0[0]\, B => 
        defSlaveSMNextState_m_0_3, C => \d_count_i_1[0]\, D => 
        d_m2_e_1, Y => \d_count_i_2[0]\);
    
    \mask[7]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(7), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[7]_net_1\);
    
    \ins2[25]\ : SLE
      port map(D => \d_ins2[25]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[25]_net_1\);
    
    \state_ns_0_0[8]\ : CFG4
      generic map(INIT => x"02F2")

      port map(A => \state[20]_net_1\, B => \state[15]_net_1\, C
         => \state[16]_net_1\, D => N_125, Y => 
        \state_ns_0_0[8]_net_1\);
    
    \haddr_fetch_RNO[8]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_6_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[8]\, D => N_4812, Y => N_4365_i_0);
    
    \haddr_fetch_RNO[14]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_s_12_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[14]\, D => N_4812, Y => 
        N_2651_i_0);
    
    \state[14]\ : SLE
      port map(D => N_16_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[14]_net_1\);
    
    \rdata[6]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(6), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[6]_net_1\);
    
    \state_RNI8H011[22]\ : CFG4
      generic map(INIT => x"4044")

      port map(A => \count[1]_net_1\, B => \state[22]_net_1\, C
         => N_4917, D => N_249, Y => N_579);
    
    \HWDATA_int_RNO_1[5]\ : CFG4
      generic map(INIT => x"8F88")

      port map(A => \state[10]_net_1\, B => \acc[5]_net_1\, C => 
        N_274, D => N_4539, Y => d_HWDATA_0_iv_25_605_7_0);
    
    un7_hready_2_RNIJCHN : CFG4
      generic map(INIT => x"4000")

      port map(A => \ins1[20]_net_1\, B => \ins1[21]_net_1\, C
         => un9_hready_2, D => \state[22]_net_1\, Y => N_403);
    
    \d_HADDR_0_iv[11]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_2[11]_net_1\, B => 
        un46_d_haddr_cry_11_S, C => \d_HADDR_0_iv_1[11]_net_1\, D
         => N_247, Y => \d_HADDR[11]\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o2 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => N_4901, B => N_252, C => N_4902, D => 
        \un1_d_HWRITE_1_sqmuxa_2_i_o2_1\, Y => N_247);
    
    \HSIZE_int_RNO[1]\ : CFG1
      generic map(INIT => "01")

      port map(A => \un7_iv_0_a1_0[14]_net_1\, Y => 
        \un7_iv_0_a1_0_i[14]\);
    
    \HADDR_int[24]\ : SLE
      port map(D => \d_HADDR[24]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[24]\);
    
    state_21_rep1_RNI8UPFA : CFG4
      generic map(INIT => x"FFEA")

      port map(A => N_290, B => \state_21_rep1\, C => 
        defSlaveSMNextState_m_0_2, D => un1_state_31_i_i_o2_0, Y
         => un1_state_31_i_i_a2_0_d_1_sx_0);
    
    un1_state_42_0_0_3 : CFG4
      generic map(INIT => x"AEFF")

      port map(A => \un1_state_42_0_0_1\, B => N_136, C => 
        HREADY_i_3, D => N_228, Y => \un1_state_42_0_0_3\);
    
    \state_RNO[7]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \state[25]_net_1\, B => \state[7]_net_1\, C
         => N_379, D => HREADY_i_3, Y => N_20_i_0);
    
    \d_HADDR_0_iv_0_0_a2[24]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[24]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_481);
    
    \state_RNIG0L12[21]\ : CFG4
      generic map(INIT => x"37FF")

      port map(A => N_252, B => N_390, C => \state[21]_net_1\, D
         => N_251, Y => d_HWDATA_0_iv_8_1298_1_o2_i_1);
    
    \state_RNIANFH[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => \state[4]_net_1\, Y => 
        N_696_i_0);
    
    \count_RNO_5[1]\ : CFG4
      generic map(INIT => x"5155")

      port map(A => N_319, B => N_259, C => N_375, D => 
        d_m2_e_2_2, Y => \d_count_0_o2_0_1_2[1]\);
    
    un1_hready_2_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \count[1]_net_1\, B => \count[0]_net_1\, Y
         => N_4912);
    
    \d_acc_1_0[16]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[16]_net_1\, B => \acc[16]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[16]_net_1\);
    
    \d_ins2[29]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(29), B => un28_opcode, 
        Y => \d_ins2[29]_net_1\);
    
    \d_acc_0[19]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[19]_net_1\, B => \ins2[19]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(19), D => \state[8]_net_1\, Y => 
        N_1156);
    
    \rdata_RNIMC2I[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \rdata[17]_net_1\, B => \count[1]_net_1\, C
         => \rdata[1]_net_1\, Y => N_388);
    
    \HWDATA_int_RNO_0[7]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_270, C => 
        \acc[7]_net_1\, D => \rdata[7]_net_1\, Y => 
        d_HWDATA_0_iv_23_695_0_0);
    
    \HWDATA_int_RNO[14]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_16_956_0_0, B => N_680_2, C => 
        \rdata[14]_net_1\, D => N_264, Y => 
        \HWDATA_int_RNO[14]_net_1\);
    
    \HADDR_int[23]\ : SLE
      port map(D => \d_HADDR[23]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[23]\);
    
    \bytecount_RNO[8]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4337, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_42_i_0);
    
    \HWDATA_int[13]\ : SLE
      port map(D => \HWDATA_int_RNO[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(13));
    
    \haddr_fetch[28]\ : SLE
      port map(D => N_19_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[28]_net_1\);
    
    \count_RNIOM5RC[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_252, B => defSlaveSMNextState_m_0_3, C => 
        \count[1]_net_1\, Y => d_m2_e_2_0_1);
    
    un1_state_44_0_8 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[6]_net_1\, B => \state[17]_net_1\, C
         => \un1_state_44_0_6\, D => \state[10]_net_1\, Y => 
        \un1_state_44_0_8\);
    
    \haddr_write[9]\ : SLE
      port map(D => un46_d_haddr_cry_9_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[9]_net_1\);
    
    \rdata_RNIPG3I[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \rdata[23]_net_1\, B => \count[1]_net_1\, C
         => \rdata[7]_net_1\, Y => N_2570);
    
    \ins1[16]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(16), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[16]_net_1\);
    
    d_bytecount_0_sqmuxa_i_o2 : CFG3
      generic map(INIT => x"DF")

      port map(A => \state[25]_net_1\, B => \ins1[25]_net_1\, C
         => N_198, Y => N_78);
    
    \HWDATA_int_RNO[7]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_23_695_0_0, B => N_285, C => 
        \rdata[23]_net_1\, D => N_271, Y => 
        \HWDATA_int_RNO[7]_net_1\);
    
    \ins1[6]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(6), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[6]_net_1\);
    
    \HWDATA_int_RNO[24]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => d_HWDATA_0_iv_6_1388_5_0, B => 
        \rdata[24]_net_1\, C => N_682_2, D => N_277, Y => N_2351);
    
    un13_d_haddr_1_cry_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[17]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_14\, S => un13_d_haddr_1_cry_15_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_15\);
    
    \state_ns[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \state[13]_net_1\, B => \state[12]_net_1\, C
         => HREADY_i_3, Y => \state_ns[16]_net_1\);
    
    un46_d_haddr_cry_20 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[20]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_19\, S => un46_d_haddr_cry_20_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_20\);
    
    \mask[3]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(3), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[3]_net_1\);
    
    \d_HADDR_0_iv_0[11]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => un13_d_haddr_1_cry_9_S, B => \state_ns[0]\, C
         => N_4814, D => \un1_state_30_0_0\, Y => 
        \d_HADDR_0_iv_0[11]_net_1\);
    
    \d_acc_1[21]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[21]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(21), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[21]\);
    
    \haddr_fetch_RNO[10]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_8_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[10]\, D => N_4812, Y => 
        N_4364_i_0);
    
    \HWDATA_int_RNO_1[0]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => \rdata[16]_net_1\, B => \rdata[0]_net_1\, C
         => N_4890, D => N_4687, Y => d_HWDATA_0_iv_30_380_1_2);
    
    un1_rdata_0_I_1 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[1]_net_1\, B => N_83_i, C => 
        \expected[1]_net_1\, D => \mask[1]_net_1\, FCI => 
        VCC_net_1, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[0]\);
    
    \d_ins2[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(3), B => un28_opcode, 
        Y => \d_ins2[3]_net_1\);
    
    \d_acc[6]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1143, C => 
        \ins2[6]_net_1\, D => \acc[6]_net_1\, Y => 
        \d_acc[6]_net_1\);
    
    \count_RNIUH5O_0[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4879, B => N_251, Y => N_4777_1);
    
    un1_rdata_0_I_70 : CFG3
      generic map(INIT => x"6A")

      port map(A => \expected[31]_net_1\, B => \rdata[31]_net_1\, 
        C => \mask[31]_net_1\, Y => un1_rdata_0_N_22);
    
    \haddr_write[20]\ : SLE
      port map(D => un46_d_haddr_cry_20_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[20]_net_1\);
    
    \rdata[25]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(25), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[25]_net_1\);
    
    \d_HADDR_0_iv_2[23]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_23_S, B => 
        \d_HADDR_0_iv_0[23]_net_1\, C => \ins2_m[23]\, D => N_247, 
        Y => \d_HADDR_0_iv_2[23]_net_1\);
    
    \d_ins2[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(5), B => un28_opcode, 
        Y => \d_ins2[5]_net_1\);
    
    \HWDATA_int_RNO_0[14]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[14]_net_1\, D => \rdata[30]_net_1\, Y => 
        d_HWDATA_0_iv_16_956_0_0);
    
    \mask[6]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(6), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[6]_net_1\);
    
    \ins1_RNI6O3UF5[7]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[7]_net_1\, B => N_78, C => N_164, 
        D => \ins1[7]_net_1\, FCI => d_bytecount_i_m2_cry_6, S
         => N_108, Y => OPEN, FCO => d_bytecount_i_m2_cry_7);
    
    \d_ins2[18]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(18), B => un28_opcode, 
        Y => \d_ins2[18]_net_1\);
    
    \haddr_write[17]\ : SLE
      port map(D => un46_d_haddr_cry_17_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[17]_net_1\);
    
    \acc[24]\ : SLE
      port map(D => \d_acc[24]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[24]_net_1\);
    
    \d_HADDR_0_iv_2_RNO[23]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[23]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[23]\);
    
    un13_d_haddr_1_cry_18 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[20]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_17\, S => un13_d_haddr_1_cry_18_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_18\);
    
    \rdata[14]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(14), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[14]_net_1\);
    
    \mask[21]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(21), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[21]_net_1\);
    
    \haddr_write[30]\ : SLE
      port map(D => un46_d_haddr_cry_30_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[30]_net_1\);
    
    \expected[19]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(19), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[19]_net_1\);
    
    un1_state_39_1_0_a3_3_0_o2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \ins1[30]_net_1\, B => \ins1[29]_net_1\, C
         => \ins1[28]_net_1\, D => \ins1[27]_net_1\, Y => N_80);
    
    \rdata_RNID9Q62[12]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \rdata[28]_net_1\, B => \rdata[12]_net_1\, C
         => N_655, D => N_600, Y => N_287);
    
    \bytecount[6]\ : SLE
      port map(D => N_38_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[6]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ins1_RNINVMUA9[12]\ : ARI1
      generic map(INIT => x"5D872")

      port map(A => \bytecount[12]_net_1\, B => N_78, C => N_164, 
        D => \ins1[12]_net_1\, FCI => d_bytecount_i_m2_cry_11, S
         => N_114, Y => OPEN, FCO => d_bytecount_i_m2_cry_12);
    
    \HADDR_int_RNO[16]\ : CFG3
      generic map(INIT => x"31")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[16]_net_1\, C => 
        \haddr_fetch[16]_net_1\, Y => \d_HADDR_0_iv_i_0[16]\);
    
    \d_HADDR_0_iv_0_0_a3_0_0[24]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \state[23]_net_1\, B => 
        \haddr_write[24]_net_1\, Y => 
        \d_HADDR_0_iv_0_0_a3_0_0[24]_net_1\);
    
    \count_RNIU5932[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_258, B => d_HWDATA_0_iv_7_1343_o2_0_0, C
         => \count[1]_net_1\, Y => N_283);
    
    \rdata_RNIMBUS1[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[19]_net_1\, B => \rdata[3]_net_1\, C
         => N_592, D => N_254, Y => N_683_2);
    
    \rdata[13]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(13), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[13]_net_1\);
    
    \d_HADDR_0_iv_0_a6_1[18]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[18]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4387);
    
    \state_RNIDD3I[22]\ : CFG4
      generic map(INIT => x"038B")

      port map(A => \state[22]_net_1\, B => \count[1]_net_1\, C
         => N_252, D => N_249, Y => \d_count_0_o3_3_0[1]\);
    
    \mask[12]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(12), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[12]_net_1\);
    
    \haddr_write[2]\ : SLE
      port map(D => un46_d_haddr_cry_2_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[2]_net_1\);
    
    \count_RNO_6[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_252, B => N_294, C => N_266, Y => N_444);
    
    \rdata[22]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(22), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[22]_net_1\);
    
    \HWDATA_int[5]\ : SLE
      port map(D => \HWDATA_int_RNO[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(5));
    
    un1_d_HWRITE_0_sqmuxa_5_i_0_0 : CFG4
      generic map(INIT => x"BA30")

      port map(A => un1_d_HWRITE_0_sqmuxa_5_i_a3_0, B => 
        HREADY_i_3, C => N_137, D => d_HWRITE_0_sqmuxa_4, Y => 
        \un1_d_HWRITE_0_sqmuxa_5_i_0_0\);
    
    \haddr_fetch[5]\ : SLE
      port map(D => \haddr_fetch_RNO[5]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[5]_net_1\);
    
    \d_bytecount[15]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_1116, B => \state[21]_net_1\, C => N_109_i, 
        Y => \d_bytecount[15]_net_1\);
    
    \rdata_RNIQJ511[30]\ : CFG4
      generic map(INIT => x"AC0F")

      port map(A => \rdata[22]_net_1\, B => \rdata[30]_net_1\, C
         => d_HWDATA_0_iv_8_1298_1_o2_i_m2_ns_1, D => 
        \count[1]_net_1\, Y => N_390);
    
    \haddr_fetch[0]\ : SLE
      port map(D => \ConfigMaster_0_M_HADDR[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[0]_net_1\);
    
    \acc[0]\ : SLE
      port map(D => \d_acc[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[0]_net_1\);
    
    \HADDR_int_RNO_0[30]\ : CFG4
      generic map(INIT => x"4445")

      port map(A => \d_HADDR_0_iv_0_0[30]_net_1\, B => 
        \haddr_fetch[30]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => \d_HADDR_0_iv_i_1[30]\);
    
    un1_d_HWRITE_0_sqmuxa_1_0_a3_i : CFG4
      generic map(INIT => x"FFFE")

      port map(A => defSlaveSMNextState_m_0_2, B => 
        defSlaveSMNextState_m_0_3, C => 
        \un1_d_HWRITE_0_sqmuxa_1_0_a3_i_1\, D => 
        un1_state_31_i_i_a2_0_d_1_0_1, Y => N_228);
    
    state_m3_i_2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \state[6]_net_1\, B => \state[27]_net_1\, C
         => \state[1]_net_1\, Y => \state_m3_i_2\);
    
    \d_acc[25]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1162, C => 
        \ins2[25]_net_1\, D => \acc[25]_net_1\, Y => 
        \d_acc[25]_net_1\);
    
    \state_ns_i_a2_13_0_a3[1]\ : CFG4
      generic map(INIT => x"0C8C")

      port map(A => d_state61_li, B => 
        \state_ns_i_a2_13_0_a3_8[1]_net_1\, C => 
        \state[16]_net_1\, D => \ins1[31]_net_1\, Y => N_917);
    
    \state_ns_i_0_a2_3_d_0[1]\ : CFG3
      generic map(INIT => x"5D")

      port map(A => N_156, B => N_117, C => 
        \state_ns_i_a2_10_i_2[1]_net_1\, Y => 
        \state_ns_i_0_a2_3_d_0[1]_net_1\);
    
    \HWDATA_int_RNO_0[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[29]_net_1\, B => \rdata[13]_net_1\, C
         => N_278, D => N_277, Y => d_HWDATA_0_iv_1_1568_0_1);
    
    \state_ns_0_a3_2_2[8]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \state[11]_net_1\, B => \state[13]_net_1\, C
         => \state[3]_net_1\, Y => \state_ns_0_a3_2_2[8]_net_1\);
    
    un1_rdata_0_I_15 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[27]_net_1\, B => N_331_i, C => 
        \expected[27]_net_1\, D => \mask[27]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[12]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[13]\);
    
    \count_RNIHAJ4[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_249, B => \count[1]_net_1\, Y => 
        \d_count_0_a3_13_0[1]\);
    
    un4_bytecount_0_o2_i_a2_RNICAG9O : CFG4
      generic map(INIT => x"222A")

      port map(A => \state[21]_net_1\, B => N_109_i, C => 
        defSlaveSMNextState_m, D => un1_state_31_i_i_a2_0_d_1_0_1, 
        Y => N_156);
    
    \HWDATA_int_RNO[16]\ : CFG4
      generic map(INIT => x"F8FF")

      port map(A => N_4625, B => \rdata[16]_net_1\, C => 
        d_HWDATA_0_iv_14_1028_3_1, D => N_178, Y => 
        \HWDATA_int_RNO[16]_net_1\);
    
    \ins1[25]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(25), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[25]_net_1\);
    
    \haddr_fetch[26]\ : SLE
      port map(D => N_21_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[26]_net_1\);
    
    \expected[27]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(27), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[27]_net_1\);
    
    un46_d_haddr_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[9]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_8\, S => un46_d_haddr_cry_9_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_9\);
    
    \d_acc_1_0[0]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[0]_net_1\, B => \acc[0]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[0]_net_1\);
    
    \mask[20]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(20), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[20]_net_1\);
    
    \HWDATA_int_RNO[8]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_22_740_6_0, B => N_682_2, C => 
        \rdata[8]_net_1\, D => N_264, Y => 
        \HWDATA_int_RNO[8]_net_1\);
    
    \state_RNO[25]\ : CFG3
      generic map(INIT => x"4A")

      port map(A => \state[26]_net_1\, B => \state[25]_net_1\, C
         => HREADY_i_3, Y => N_70_i_0);
    
    state_m2_e_0 : CFG3
      generic map(INIT => x"02")

      port map(A => \ins1[26]_net_1\, B => \ins1[25]_net_1\, C
         => N_80, Y => \state_m2_e_0\);
    
    HWRITE_int : SLE
      port map(D => N_727_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_31, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        ConfigMaster_0_M_HWRITE);
    
    \d_HADDR_0_iv_0[26]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_24_S, B => 
        \haddr_write[26]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[26]_net_1\);
    
    \HWDATA_int_RNO[26]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \rdata[26]_net_1\, B => N_4777_1, C => 
        d_HWDATA_0_iv_4_1460_5_2, D => N_4556_1, Y => 
        \HWDATA_int_RNO[26]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_5_i_a3_1_0 : CFG2
      generic map(INIT => x"8")

      port map(A => N_276, B => \count[1]_net_1\, Y => 
        \un1_d_HWRITE_0_sqmuxa_5_i_a3_1_0\);
    
    \HSIZE_int[1]\ : SLE
      port map(D => \un7_iv_0_a1_0_i[14]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_34_0_0\, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HSIZE(1));
    
    \d_HADDR_0_iv_0_2[16]\ : CFG4
      generic map(INIT => x"FCFD")

      port map(A => un46_d_haddr_cry_16_S, B => 
        \d_HADDR_0_iv_0_0[16]_net_1\, C => N_4759, D => N_247, Y
         => \d_HADDR_0_iv_0_2[16]_net_1\);
    
    un1_rdata_0_I_26_i_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[15]_net_1\, B => \rdata[15]_net_1\, 
        C => \mask[15]_net_1\, Y => N_339_i);
    
    \state_RNIPNVM[22]\ : CFG3
      generic map(INIT => x"D5")

      port map(A => \state[22]_net_1\, B => \state[21]_net_1\, C
         => N_249, Y => N_281);
    
    \d_ins2[24]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(24), B => un28_opcode, 
        Y => \d_ins2[24]_net_1\);
    
    \d_HADDR_0_iv_0[28]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_26_S, B => 
        \haddr_write[28]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0[28]_net_1\);
    
    \state_ns_0_0_a2_0_2[17]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \ins1[25]_net_1\, B => \ins1[26]_net_1\, C
         => N_654, D => N_80, Y => N_411_2);
    
    \d_acc_0[26]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[26]_net_1\, B => \ins2[26]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(26), D => \state[8]_net_1\, Y => 
        N_1163);
    
    un1_state_25_0_0 : CFG3
      generic map(INIT => x"CE")

      port map(A => \state[12]_net_1\, B => N_789, C => 
        HREADY_i_3, Y => \un1_state_25_0_0\);
    
    \d_acc_1_a2_0_0[10]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \state[7]_net_1\, B => \state[8]_net_1\, Y
         => \d_acc_1_a2_0_0[5]\);
    
    \d_acc[31]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1168, C => 
        \ins2[31]_net_1\, D => \acc[31]_net_1\, Y => 
        \d_acc[31]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_1_0 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => N_404, B => N_403, C => N_228, D => N_402, Y
         => \un1_d_HWRITE_0_sqmuxa_1_0\);
    
    \d_HADDR_0_iv_2_RNO[9]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[9]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[9]\);
    
    \count_RNIUH5O[0]\ : CFG4
      generic map(INIT => x"DDCD")

      port map(A => \state[21]_net_1\, B => \count[0]_net_1\, C
         => N_252, D => N_4711, Y => N_4890);
    
    d_count_1_sqmuxa_i_a2_0_o2_i_o2_RNIPGTI : CFG4
      generic map(INIT => x"0040")

      port map(A => \state[21]_net_1\, B => \count[0]_net_1\, C
         => N_252, D => N_259, Y => N_4917);
    
    \HWDATA_int_RNO[11]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_19_848_6_0, B => N_683_2, C => 
        \rdata[11]_net_1\, D => N_264, Y => N_1926);
    
    un1_d_HTRANS_0_sqmuxa_i_a2_0_i_o3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[12]_net_1\, B => \state[9]_net_1\, C
         => \state[7]_net_1\, D => \state[8]_net_1\, Y => N_117);
    
    \d_HADDR_0_iv_0_2[13]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[13]_net_1\, B => 
        \ins2[13]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_0_2[13]_net_1\);
    
    \d_acc_0[31]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[31]_net_1\, B => \ins2[31]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(31), D => \state[8]_net_1\, Y => 
        N_1168);
    
    \count_RNO_8[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_249, B => N_272, Y => \d_count_0_a2_2_0[1]\);
    
    \count_RNO_4[0]\ : CFG4
      generic map(INIT => x"0257")

      port map(A => \count[0]_net_1\, B => \state[21]_net_1\, C
         => N_259, D => N_542_2, Y => \d_count_i_a2_2_1_0[0]\);
    
    \d_HADDR_0_iv_2_RNO[26]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[26]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[26]\);
    
    \state_RNO[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => d_state61_li, B => \state[16]_net_1\, Y => 
        \state_ns[13]\);
    
    \state[7]\ : SLE
      port map(D => N_20_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[7]_net_1\);
    
    \rdata_RNI94ME[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \state[22]_net_1\, B => \rdata[15]_net_1\, Y
         => N_2573_1);
    
    \ins2[21]\ : SLE
      port map(D => \d_ins2[21]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[21]_net_1\);
    
    \ins2[23]\ : SLE
      port map(D => \d_ins2[23]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[23]_net_1\);
    
    \d_HADDR_0_iv_RNO[27]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => un13_d_haddr_1_cry_25_S, B => 
        \un1_state_30_0_0\, C => N_4814, Y => 
        \un13_d_haddr_1_m[27]\);
    
    \HWDATA_int_RNO[21]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_9_1253_1_1, B => N_2246_1, C
         => \rdata[21]_net_1\, D => N_403, Y => 
        \HWDATA_int_RNO[21]_net_1\);
    
    \d_HADDR_0_iv_0_0[10]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => un13_d_haddr_1_cry_8_S, B => 
        \haddr_write[10]_net_1\, C => N_4874, D => un1_state_30, 
        Y => \d_HADDR_0_iv_0_0[10]_net_1\);
    
    \d_HADDR_0_iv_0_1_0[7]\ : CFG4
      generic map(INIT => x"1115")

      port map(A => N_4592, B => \haddr_fetch[7]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => 
        \d_HADDR_0_iv_0_1_0[7]_net_1\);
    
    \ins2[28]\ : SLE
      port map(D => \d_ins2[28]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[28]_net_1\);
    
    un46_d_haddr_cry_21 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[21]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_20\, S => un46_d_haddr_cry_21_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_21\);
    
    \HWDATA_int_RNO[10]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_20_812_0_0, B => N_4556_1, C
         => \rdata[10]_net_1\, D => N_264, Y => N_1897);
    
    \count_RNO[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_453, B => N_452, C => \d_count_i_2[0]\, D
         => N_450, Y => N_4888_i_0);
    
    \d_acc_1_0[13]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[13]_net_1\, B => \acc[13]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[13]_net_1\);
    
    \rdata[21]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(21), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[21]_net_1\);
    
    \haddr_fetch_RNO[27]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_25_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[27]\, D => N_4812, Y => 
        N_4407_i_0);
    
    \mask[19]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(19), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[19]_net_1\);
    
    \rdata_RNIG5US1[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[16]_net_1\, B => \rdata[0]_net_1\, C
         => N_592, D => N_254, Y => N_682_2);
    
    \HADDR_int[26]\ : SLE
      port map(D => \d_HADDR[26]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[26]\);
    
    \count_RNIQKL51[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_255, B => \count[1]_net_1\, Y => N_601);
    
    \HWDATA_int_RNO[20]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \rdata[4]_net_1\, B => N_601, C => 
        d_HWDATA_0_iv_10_1208_0_1, D => N_287, Y => 
        \HWDATA_int_RNO[20]_net_1\);
    
    \expected[10]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(10), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[10]_net_1\);
    
    \d_HADDR_0_iv_0_2[17]\ : CFG4
      generic map(INIT => x"FCFD")

      port map(A => un46_d_haddr_cry_17_S, B => 
        \d_HADDR_0_iv_0_0[17]_net_1\, C => \ins2_i_m[17]\, D => 
        N_247, Y => \d_HADDR_0_iv_0_2[17]_net_1\);
    
    \state_RNI9MFH[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => HREADY_i_3, B => \state[3]_net_1\, Y => 
        N_14_i_0);
    
    \ins2[15]\ : SLE
      port map(D => \d_ins2[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[15]_net_1\);
    
    \HWDATA_int[0]\ : SLE
      port map(D => \HWDATA_int_RNO[0]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(0));
    
    \rdata[4]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(4), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[4]_net_1\);
    
    \HWDATA_int_RNO_0[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[11]_net_1\, D => \rdata[27]_net_1\, Y => 
        d_HWDATA_0_iv_19_848_6_0);
    
    \bytecount_RNO[6]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_4336, B => \state[21]_net_1\, C => N_109_i, 
        Y => N_38_i_0);
    
    \state[11]\ : SLE
      port map(D => \state_ns[17]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[11]_net_1\);
    
    \pause_count[3]\ : SLE
      port map(D => N_4808_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        pause_counte, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pause_count[3]_net_1\);
    
    \HADDR_int[3]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[3]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[3]\);
    
    \d_HADDR_0_iv_1[15]\ : CFG4
      generic map(INIT => x"0357")

      port map(A => \haddr_write[15]_net_1\, B => 
        \ins2[15]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_1[15]_net_1\);
    
    \HWDATA_int_RNO_0[17]\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => N_512_1, B => N_4625, C => \rdata[17]_net_1\, 
        D => N_475, Y => d_HWDATA_0_iv_13_1073_0_1);
    
    \HADDR_int[31]\ : SLE
      port map(D => \d_HADDR[31]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[31]\);
    
    \d_acc[8]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1145, C => 
        \ins2[8]_net_1\, D => \acc[8]_net_1\, Y => 
        \d_acc[8]_net_1\);
    
    \expected[29]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(29), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[29]_net_1\);
    
    \HWDATA_int_RNO_0[24]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_278, C => 
        \acc[24]_net_1\, D => \rdata[8]_net_1\, Y => 
        d_HWDATA_0_iv_6_1388_5_0);
    
    \d_acc_1_0[30]\ : CFG4
      generic map(INIT => x"EE80")

      port map(A => \ins2[30]_net_1\, B => \acc[30]_net_1\, C => 
        \state[8]_net_1\, D => \state[7]_net_1\, Y => 
        \d_acc_1_0[30]_net_1\);
    
    \count_RNITHHQA[0]\ : CFG3
      generic map(INIT => x"04")

      port map(A => un1_state_31_i_i_a2_0_d_1_0_1, B => 
        \count[0]_net_1\, C => defSlaveSMNextState_m_0_2, Y => 
        d_m2_e_1);
    
    \acc[12]\ : SLE
      port map(D => \d_acc[12]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[12]_net_1\);
    
    \d_ins2[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(28), B => un28_opcode, 
        Y => \d_ins2[28]_net_1\);
    
    \state_ns_i_a2_13_0_a3_5_0[1]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \state[3]_net_1\, B => \state[19]_net_1\, C
         => \state[17]_net_1\, D => \state[15]_net_1\, Y => 
        \state_ns_i_a2_13_0_a3_5_0[1]_net_1\);
    
    \rdata_RNIA7R62[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[31]_net_1\, B => \rdata[15]_net_1\, C
         => N_600, D => N_655, Y => N_285);
    
    \HADDR_int_RNO_0[6]\ : CFG4
      generic map(INIT => x"4445")

      port map(A => \d_HADDR_0_iv_0[6]_net_1\, B => 
        \haddr_fetch[6]_net_1\, C => 
        \un1_d_HWRITE_0_sqmuxa_2_0_0\, D => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, Y => \d_HADDR_0_iv_i_1[6]\);
    
    un46_d_haddr_cry_3_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[19]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[3]\, C => GND_net_1, D => 
        GND_net_1, FCI => un46_d_haddr_cry_2_0_FCO, S => OPEN, Y
         => OPEN, FCO => un46_d_haddr_cry_3_0_FCO);
    
    \HTRANS_int[1]\ : SLE
      port map(D => \un1_state_42_0_0\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_46\, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ConfigMaster_0_M_HTRANS(1));
    
    un1_state_44_0_4 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[28]_net_1\, B => \state[20]_net_1\, C
         => \state[15]_net_1\, D => \state[3]_net_1\, Y => 
        \un1_state_44_0_4\);
    
    un1_d_haddr_fetch_2_sqmuxa : CFG4
      generic map(INIT => x"0EFF")

      port map(A => \d_haddr_fetch_2_sqmuxa_0\, B => N_4812, C
         => HREADY_i_3, D => N_78, Y => 
        \un1_d_haddr_fetch_2_sqmuxa\);
    
    \d_HADDR_0_iv_0_2[5]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => un46_d_haddr_cry_5_S, B => 
        \d_HADDR_0_iv_0_0[5]_net_1\, C => N_4524, D => N_247, Y
         => \d_HADDR_0_iv_0_2[5]_net_1\);
    
    un1_state_44_0_6 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \state[13]_net_1\, B => \state[18]_net_1\, C
         => \state[2]_net_1\, D => \state[4]_net_1\, Y => 
        \un1_state_44_0_6\);
    
    un46_d_haddr_cry_17 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[17]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_16\, S => un46_d_haddr_cry_17_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_17\);
    
    un1_state_34_0_a2_0_0_a3 : CFG4
      generic map(INIT => x"0200")

      port map(A => \state[21]_net_1\, B => \ins1[31]_net_1\, C
         => HREADY_i_3, D => N_109_i, Y => N_929);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o3_1_1 : CFG3
      generic map(INIT => x"A2")

      port map(A => \count[1]_net_1\, B => N_249, C => 
        \count[0]_net_1\, Y => un1_d_HWRITE_1_sqmuxa_2_i_o3_1_0);
    
    un46_d_haddr_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[13]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_12\, S => un46_d_haddr_cry_13_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_13\);
    
    \state_ns_a2_1_i_o2_0[4]\ : CFG4
      generic map(INIT => x"555D")

      port map(A => \state[25]_net_1\, B => \ins1[26]_net_1\, C
         => N_80, D => \ins1[25]_net_1\, Y => N_86);
    
    \rdata_RNIR9Q5[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \count[1]_net_1\, B => \rdata[21]_net_1\, Y
         => N_4541);
    
    \HWDATA_int_RNO_0[30]\ : CFG4
      generic map(INIT => x"B3A0")

      port map(A => \state[10]_net_1\, B => N_263, C => 
        \acc[30]_net_1\, D => \rdata[14]_net_1\, Y => 
        d_HWDATA_0_iv_0_1604_5_0);
    
    \expected[14]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(14), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[14]_net_1\);
    
    un1_d_HWRITE_0_sqmuxa_5_i_a3_0_0 : CFG4
      generic map(INIT => x"1113")

      port map(A => \state[21]_net_1\, B => \state[10]_net_1\, C
         => d_state_1_sqmuxa_1_i_0, D => N_109_i, Y => 
        un1_d_HWRITE_0_sqmuxa_5_i_a3_0);
    
    d_HWRITE_0_sqmuxa_4_0_a2_1 : CFG4
      generic map(INIT => x"0080")

      port map(A => N_661, B => \state[22]_net_1\, C => 
        d_N_3_mux_0, D => N_249, Y => N_404);
    
    \expected[16]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(16), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[16]_net_1\);
    
    \d_HADDR_0_iv[2]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[2]_net_1\, C => \haddr_fetch[2]_net_1\, Y
         => \d_HADDR[2]\);
    
    \HADDR_int[25]\ : SLE
      port map(D => \d_HADDR[25]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[25]\);
    
    un46_d_haddr_cry_18 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[18]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_17\, S => un46_d_haddr_cry_18_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_18\);
    
    \haddr_fetch[2]\ : SLE
      port map(D => N_64_i, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[2]_net_1\);
    
    \haddr_fetch[7]\ : SLE
      port map(D => \haddr_fetch_RNO[7]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[7]_net_1\);
    
    \haddr_fetch[19]\ : SLE
      port map(D => N_4367_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[19]_net_1\);
    
    \rdata[3]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(3), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[3]_net_1\);
    
    \HADDR_int[14]\ : SLE
      port map(D => \d_HADDR[14]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[14]\);
    
    \bytecount[3]\ : SLE
      port map(D => \d_bytecount[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[3]_net_1\);
    
    \pause_count[1]\ : SLE
      port map(D => N_37_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        pause_counte, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pause_count[1]_net_1\);
    
    \HWDATA_int[27]\ : SLE
      port map(D => \HWDATA_int_RNO[27]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(27));
    
    \d_ins2[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(10), B => un28_opcode, 
        Y => \d_ins2[10]_net_1\);
    
    \ins1[21]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(21), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[21]_net_1\);
    
    \state_ns_0[7]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \state[21]_net_1\, B => 
        d_state_1_sqmuxa_1_i_0, C => N_109_i, D => N_101, Y => 
        \state_ns[7]\);
    
    \ins2[27]\ : SLE
      port map(D => \d_ins2[27]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[27]_net_1\);
    
    \HWDATA_int[4]\ : SLE
      port map(D => \HWDATA_int_RNO[4]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(4));
    
    \ins1[23]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(23), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[23]_net_1\);
    
    \haddr_fetch_RNO[18]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_16_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[18]\, D => N_4812, Y => 
        \haddr_fetch_RNO[18]_net_1\);
    
    \acc[6]\ : SLE
      port map(D => \d_acc[6]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[6]_net_1\);
    
    \HADDR_int[13]\ : SLE
      port map(D => \d_HADDR[13]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[13]\);
    
    \d_HADDR_0_iv_0_a2_3[21]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[21]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4514);
    
    \HWDATA_int_RNO[9]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => N_2380_3, B => \rdata[9]_net_1\, C => 
        d_HWDATA_0_iv_21_776_6_0, D => N_264, Y => 
        \HWDATA_int_RNO[9]_net_1\);
    
    \ins1[28]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(28), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[28]_net_1\);
    
    \rdata[8]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(8), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[8]_net_1\);
    
    \state_RNI3IUI[19]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \state[19]_net_1\, B => \state[23]_net_1\, Y
         => N_4812);
    
    \ins1[2]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(2), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[2]_net_1\);
    
    \HWDATA_int_RNO[13]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => N_301, B => \rdata[13]_net_1\, C => 
        d_HWDATA_0_iv_17_920_0_0, D => N_264, Y => 
        \HWDATA_int_RNO[13]_net_1\);
    
    \d_HADDR_0_iv_0_0[0]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => \ConfigMaster_0_M_HADDR[0]\, B => 
        \haddr_write[0]_net_1\, C => N_4874, D => un1_state_30, Y
         => \d_HADDR_0_iv_0_0[0]_net_1\);
    
    \acc[20]\ : SLE
      port map(D => \d_acc[20]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[20]_net_1\);
    
    \rdata_RNIBK3K1[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \rdata[21]_net_1\, B => N_4472, C => N_4916, 
        D => N_656, Y => N_301);
    
    \HWDATA_int_RNO[31]\ : CFG4
      generic map(INIT => x"FFB3")

      port map(A => N_4777_1, B => d_HWDATA_0_iv_1640_1, C => 
        \rdata[31]_net_1\, D => N_2061, Y => 
        \HWDATA_int_RNO[31]_net_1\);
    
    \haddr_write[25]\ : SLE
      port map(D => un46_d_haddr_cry_25_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[25]_net_1\);
    
    \haddr_write[12]\ : SLE
      port map(D => un46_d_haddr_cry_12_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[12]_net_1\);
    
    \HWDATA_int_RNO_0[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_4687, C => 
        \acc[6]_net_1\, D => \rdata[6]_net_1\, Y => 
        d_HWDATA_0_iv_24_650_7_0);
    
    un13_d_haddr_1_cry_27 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[29]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_26\, S => un13_d_haddr_1_cry_27_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_27\);
    
    un1_rdata_0_I_20_i_0_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[26]_net_1\, B => \rdata[26]_net_1\, 
        C => \mask[26]_net_1\, Y => N_331_i);
    
    \state[27]\ : SLE
      port map(D => N_741_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[27]_net_1\);
    
    \HWDATA_int_RNO[23]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_7_1343_1_0, B => N_285, C => 
        \rdata[23]_net_1\, D => N_283, Y => 
        \HWDATA_int_RNO[23]_net_1\);
    
    \haddr_fetch_RNO[22]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_20_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[22]\, D => N_4812, Y => 
        N_4722_i_0);
    
    \count_RNIGSAG2[0]\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => N_249, B => d_HWDATA_0_iv_8_1298_1_o2_i_1, C
         => \count[0]_net_1\, D => N_263, Y => N_4891);
    
    \rdata[26]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(26), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[26]_net_1\);
    
    \d_ins2[17]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(17), B => un28_opcode, 
        Y => \d_ins2[17]_net_1\);
    
    \d_HADDR_0_iv_1[31]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[31]_net_1\, B => 
        \ins2[31]_net_1\, C => N_4873, D => N_4874, Y => 
        \d_HADDR_0_iv_1[31]_net_1\);
    
    \d_acc_1[30]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \d_acc_1_0[30]_net_1\, B => 
        ConfigMaster_0_M_HRDATA(30), C => \d_acc_1_a2_0_0[5]\, Y
         => \d_acc[30]\);
    
    un46_d_haddr_cry_2_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => \ins1[18]_net_1\, B => 
        \ConfigMaster_0_M_HADDR[2]\, C => GND_net_1, D => 
        GND_net_1, FCI => un46_d_haddr_cry_1_0_FCO, S => OPEN, Y
         => OPEN, FCO => un46_d_haddr_cry_2_0_FCO);
    
    \HWDATA_int[3]\ : SLE
      port map(D => \HWDATA_int_RNO[3]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(3));
    
    HWRITE_int_RNO : CFG3
      generic map(INIT => x"0E")

      port map(A => \state[11]_net_1\, B => N_259, C => 
        HREADY_i_3, Y => N_727_i_0);
    
    \d_acc_0[8]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[8]_net_1\, B => \ins2[8]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(8), D => \state[8]_net_1\, Y => 
        N_1145);
    
    \count_RNIQB601[1]\ : CFG4
      generic map(INIT => x"5450")

      port map(A => \count[1]_net_1\, B => \state[21]_net_1\, C
         => N_674, D => N_249, Y => N_600);
    
    un1_rdata_0_I_93 : ARI1
      generic map(INIT => x"48222")

      port map(A => \rdata[24]_net_1\, B => N_327_i, C => 
        \expected[24]_net_1\, D => \mask[24]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[11]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[12]\);
    
    \pause_count_RNO[0]\ : CFG3
      generic map(INIT => x"07")

      port map(A => N_4813, B => \pause_count[0]_net_1\, C => 
        N_3400, Y => N_4316_i_0);
    
    un1_state_46_1 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \un1_state_46_0\, B => HREADY_i_3, C => 
        \ins1[31]_net_1\, D => N_789, Y => \un1_state_46_1\);
    
    un12_size_2_0_5 : CFG4
      generic map(INIT => x"0001")

      port map(A => \bytecount[11]_net_1\, B => 
        \bytecount[10]_net_1\, C => \bytecount[9]_net_1\, D => 
        \bytecount[8]_net_1\, Y => \un12_size_2_0_5\);
    
    \HWDATA_int_RNO[30]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => d_HWDATA_0_iv_0_1604_5_0, B => N_4778, C => 
        d_HWDATA_0_iv_0_1604_1_0, D => N_680_2, Y => N_2525);
    
    \HWDATA_int[24]\ : SLE
      port map(D => N_2351, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(24));
    
    un13_d_haddr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[9]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_6\, S => un13_d_haddr_1_cry_7_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_7\);
    
    \haddr_fetch_RNO[21]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_19_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[21]\, D => N_4812, Y => N_62);
    
    \expected[20]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(20), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[20]_net_1\);
    
    \count_RNO_6[0]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => N_266, B => \state[21]_net_1\, C => N_290, D
         => N_259, Y => \d_count_i_a2_1_0[0]\);
    
    \haddr_fetch[23]\ : SLE
      port map(D => N_3216_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[23]_net_1\);
    
    \acc[29]\ : SLE
      port map(D => \d_acc[29]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[29]_net_1\);
    
    \HWDATA_int_RNO_1[30]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[22]_net_1\, B => \rdata[14]_net_1\, C
         => N_276, D => \count[1]_net_1\, Y => N_4778);
    
    \state[3]\ : SLE
      port map(D => \state[4]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        HREADY_i_3_i_0, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[3]_net_1\);
    
    \state_ns_0_a3_0[9]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ins1[25]_net_1\, B => N_198, C => N_96, D
         => HREADY_i_3, Y => N_4837);
    
    \expected[3]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(3), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[3]_net_1\);
    
    \ins1[12]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(12), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[12]_net_1\);
    
    \d_HADDR_0_iv[8]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \d_HADDR_0_iv_2[8]_net_1\, B => 
        un46_d_haddr_cry_8_S, C => \d_HADDR_0_iv_1[8]_net_1\, D
         => N_247, Y => \d_HADDR[8]\);
    
    un1_state_39_1_0_a3_1 : CFG4
      generic map(INIT => x"0200")

      port map(A => \un9_opcode_0_a2_0\, B => N_80, C => 
        \ins1[26]_net_1\, D => \state[25]_net_1\, Y => N_191);
    
    \HWDATA_int_RNO_0[21]\ : CFG4
      generic map(INIT => x"CCEC")

      port map(A => N_252, B => d_HWDATA_0_iv_9_1253_1_0, C => 
        N_4539, D => N_274, Y => d_HWDATA_0_iv_9_1253_1_1);
    
    \expected[30]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(30), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[30]_net_1\);
    
    \HWDATA_int_RNO_0[27]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_3_1496_0_0, B => N_4431, C => 
        \rdata[27]_net_1\, D => N_403, Y => 
        d_HWDATA_0_iv_3_1496_0_2);
    
    \state_RNICC3I[22]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \state[22]_net_1\, B => \count[0]_net_1\, C
         => N_252, D => N_249, Y => N_674);
    
    \HWDATA_int_RNO_0[3]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_270, C => 
        \acc[3]_net_1\, D => \rdata[3]_net_1\, Y => 
        d_HWDATA_0_iv_27_515_0_0);
    
    \haddr_fetch[21]\ : SLE
      port map(D => N_62, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[21]_net_1\);
    
    \ins2[2]\ : SLE
      port map(D => \d_ins2[2]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[2]_net_1\);
    
    \ins2[11]\ : SLE
      port map(D => \d_ins2[11]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[11]_net_1\);
    
    \haddr_fetch_RNO[29]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_27_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[29]\, D => N_4812, Y => N_18_i_0);
    
    \haddr_fetch_RNO[26]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_24_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[26]\, D => N_4812, Y => N_21_i_0);
    
    \d_ins2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(0), B => un28_opcode, 
        Y => \d_ins2[0]_net_1\);
    
    \ins2[13]\ : SLE
      port map(D => \d_ins2[13]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[13]_net_1\);
    
    state_m3_i_7 : CFG3
      generic map(INIT => x"FD")

      port map(A => N_86, B => N_4855, C => \state_m3_i_4\, Y => 
        \state_m3_i_7\);
    
    \HWDATA_int[1]\ : SLE
      port map(D => \HWDATA_int_RNO[1]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(1));
    
    busy_RNIFH7O : CFG2
      generic map(INIT => x"8")

      port map(A => \state[1]_net_1\, B => \busy\, Y => N_3400);
    
    un46_d_haddr_s_31 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[31]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_30\, S => un46_d_haddr_s_31_S, Y => 
        OPEN, FCO => OPEN);
    
    un1_d_pause_count_1_sqmuxa_i_a2_0_0_a3 : CFG4
      generic map(INIT => x"0080")

      port map(A => \state[0]_net_1\, B => \pause_count[4]_net_1\, 
        C => \pause_count[3]_net_1\, D => N_4811, Y => 
        \state_ns[22]\);
    
    \d_HADDR_0_iv_0_2[0]\ : CFG4
      generic map(INIT => x"FCFE")

      port map(A => \un46_d_haddr_axb_0\, B => 
        \d_HADDR_0_iv_0_0[0]_net_1\, C => N_4764, D => N_247, Y
         => \d_HADDR_0_iv_0_2[0]_net_1\);
    
    \ins2[18]\ : SLE
      port map(D => \d_ins2[18]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[18]_net_1\);
    
    \HWDATA_int_RNO[4]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => d_HWDATA_0_iv_26_560_0_0, B => N_287, C => 
        \rdata[20]_net_1\, D => N_271, Y => 
        \HWDATA_int_RNO[4]_net_1\);
    
    un13_d_haddr_1_s_1_172 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[2]\, 
        C => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un13_d_haddr_1_s_1_172_FCO);
    
    \HADDR_int_RNO[17]\ : CFG3
      generic map(INIT => x"31")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[17]_net_1\, C => 
        \haddr_fetch[17]_net_1\, Y => \d_HADDR_0_iv_i_0[17]\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_a2_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => N_661, B => N_249, C => d_N_3_mux_0, D => 
        N_294, Y => N_4902);
    
    \rdata[9]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(9), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[9]_net_1\);
    
    \expected[24]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(24), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[24]_net_1\);
    
    \ins1[14]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(14), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[14]_net_1\);
    
    \expected[26]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(26), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[26]_net_1\);
    
    d_count_1_sqmuxa_i_a2_0_o2_i_o2_RNIG2122 : CFG4
      generic map(INIT => x"CCEC")

      port map(A => N_291, B => N_579, C => \count[1]_net_1\, D
         => N_259, Y => \d_count_0_o2_0[1]\);
    
    \d_acc_1[16]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_789, B => \d_acc_1_0[16]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(16), Y => \d_acc[16]\);
    
    \d_acc[20]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1157, C => 
        \ins2[20]_net_1\, D => \acc[20]_net_1\, Y => 
        \d_acc[20]_net_1\);
    
    \haddr_fetch_RNO[30]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_28_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[30]\, D => N_4812, Y => N_17_i_0);
    
    \HWDATA_int_RNO_0[12]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \state[10]_net_1\, B => N_587, C => 
        \acc[12]_net_1\, D => \rdata[28]_net_1\, Y => 
        d_HWDATA_0_iv_18_884_6_0);
    
    un1_rdata_0_I_51 : ARI1
      generic map(INIT => x"40095")

      port map(A => un1_rdata_0_N_37, B => \expected[8]_net_1\, C
         => \mask[8]_net_1\, D => \rdata[8]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[3]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[4]\);
    
    \HWDATA_int_RNO_1[16]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \rdata[0]_net_1\, B => \count[1]_net_1\, C
         => N_274, D => N_252, Y => N_4741);
    
    \haddr_fetch[20]\ : SLE
      port map(D => N_4560_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[20]_net_1\);
    
    \d_HADDR_0_iv_0_a2_3[5]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[5]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => N_4524);
    
    un1_rdata_0_I_14_i_0_x2 : CFG3
      generic map(INIT => x"95")

      port map(A => \expected[28]_net_1\, B => \rdata[28]_net_1\, 
        C => \mask[28]_net_1\, Y => N_355_i);
    
    \d_HADDR_0_iv_0[12]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_0_2[12]_net_1\, C => 
        \haddr_fetch[12]_net_1\, Y => \d_HADDR[12]\);
    
    un1_d_HWRITE_0_sqmuxa_5_i_0 : CFG4
      generic map(INIT => x"FFF4")

      port map(A => HREADY_i_3, B => \state_ns_0_a2_0_1[5]_net_1\, 
        C => \un1_d_HWRITE_0_sqmuxa_5_i_0_2\, D => 
        \un1_d_HWRITE_0_sqmuxa_5_i_0_0\, Y => N_31);
    
    \mask[5]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(5), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[5]_net_1\);
    
    un46_d_haddr_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[12]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_11\, S => un46_d_haddr_cry_12_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_12\);
    
    \rdata[10]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(10), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[10]_net_1\);
    
    \mask[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[0]_net_1\);
    
    \ins1[27]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(27), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[27]_net_1\);
    
    \HWDATA_int[12]\ : SLE
      port map(D => \HWDATA_int_RNO[12]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(12));
    
    un1_rdata_0_I_81 : ARI1
      generic map(INIT => x"40095")

      port map(A => un1_rdata_0_N_12, B => \expected[4]_net_1\, C
         => \mask[4]_net_1\, D => \rdata[4]_net_1\, FCI => 
        \un1_rdata_0_data_tmp[1]\, S => OPEN, Y => OPEN, FCO => 
        \un1_rdata_0_data_tmp[2]\);
    
    \mask[23]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(23), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[23]_net_1\);
    
    \haddr_fetch_RNO[15]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_13_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[15]\, D => N_4812, Y => 
        N_4342_i_0);
    
    \state_ns_0_a3_2[8]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \state_ns_0_a3_2_2[8]_net_1\, B => 
        \state_ns_0_a3_2_3[8]_net_1\, C => N_200, D => N_212, Y
         => N_186);
    
    \mask[28]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(28), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[28]_net_1\);
    
    \count_RNI96OF1[0]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \state[21]_net_1\, B => \count[0]_net_1\, C
         => N_255, D => \count[1]_net_1\, Y => N_271);
    
    \bytecount_RNO[0]\ : CFG3
      generic map(INIT => x"70")

      port map(A => \state[21]_net_1\, B => N_109_i, C => 
        \ins1_RNIE4ISO_Y[0]\, Y => N_28_i_0);
    
    \d_HADDR_0_iv_2_RNO[25]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \ins2[25]_net_1\, B => N_837, C => HREADY_i_3, 
        Y => \ins2_m[25]\);
    
    un1_d_HWRITE_1_sqmuxa_2_i_o3_0 : CFG2
      generic map(INIT => x"B")

      port map(A => N_263, B => \count[0]_net_1\, Y => 
        \un1_d_HWRITE_1_sqmuxa_2_i_o3_0\);
    
    un9_opcode_0_a2_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \ins1[25]_net_1\, B => \ins1[24]_net_1\, Y
         => \un9_opcode_0_a2_0\);
    
    un1_state_44_0_10 : CFG4
      generic map(INIT => x"FCDC")

      port map(A => d_state61_li, B => \un1_state_44_0_9\, C => 
        \state[16]_net_1\, D => \ins1[31]_net_1\, Y => 
        \un1_state_44_0_10\);
    
    \d_acc_0[29]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => \acc[29]_net_1\, B => \ins2[29]_net_1\, C => 
        ConfigMaster_0_M_HRDATA(29), D => \state[8]_net_1\, Y => 
        N_1166);
    
    \expected[15]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(15), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[15]_net_1\);
    
    \expected[0]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(0), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[0]_net_1\);
    
    \state_RNIGI2A[22]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \count[0]_net_1\, B => \state[22]_net_1\, Y
         => N_274);
    
    \pause_count[2]\ : SLE
      port map(D => N_4807_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        pause_counte, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pause_count[2]_net_1\);
    
    \HWDATA_int[26]\ : SLE
      port map(D => \HWDATA_int_RNO[26]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(26));
    
    \mask[2]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(2), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_167, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \mask[2]_net_1\);
    
    \expected[2]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(2), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \expected[2]_net_1\);
    
    \d_acc[11]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1148, C => 
        \ins2[11]_net_1\, D => \acc[11]_net_1\, Y => 
        \d_acc[11]_net_1\);
    
    \count_RNO_5[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => N_4916, B => N_369, C => N_543, D => 
        d_N_3_mux_0, Y => \d_count_i_a2_2_1[0]\);
    
    \state_RNIP2541[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_3400, B => \state[0]_net_1\, Y => 
        pause_counte);
    
    d_HTRANS_0_sqmuxa_4_1_1_o3_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \bytecount[6]_net_1\, B => 
        \bytecount[7]_net_1\, Y => \d_HTRANS_0_sqmuxa_4_1_1_o3_1\);
    
    \state_ns_a2_0_a2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \state[1]_net_1\, B => \busy\, Y => 
        \state_ns[0]\);
    
    \ins1_RNIEV2E[22]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_274, B => N_290, Y => N_4916);
    
    \d_HADDR_0_iv[19]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[19]_net_1\, C => \haddr_fetch[19]_net_1\, 
        Y => \d_HADDR[19]\);
    
    \d_ins2[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(20), B => un28_opcode, 
        Y => \d_ins2[20]_net_1\);
    
    \d_HADDR_0_iv_1[1]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \haddr_write[1]_net_1\, B => \ins2[1]_net_1\, 
        C => N_4873, D => N_4874, Y => \d_HADDR_0_iv_1[1]_net_1\);
    
    \rdata_RNI88R71[29]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => N_4525, B => \rdata[29]_net_1\, C => N_272, Y
         => N_47);
    
    \ins1[31]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(31), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[31]_net_1\);
    
    \d_acc[27]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1164, C => 
        \ins2[27]_net_1\, D => \acc[27]_net_1\, Y => 
        \d_acc[27]_net_1\);
    
    \ins1[9]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(9), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_700_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins1[9]_net_1\);
    
    \HADDR_int[4]\ : SLE
      port map(D => \d_HADDR[4]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[4]\);
    
    \d_ins2[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(16), B => un28_opcode, 
        Y => \d_ins2[16]_net_1\);
    
    \d_HADDR_0_iv[22]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \un13_d_haddr_1_m[22]\, B => 
        un46_d_haddr_cry_22_S, C => \d_HADDR_0_iv_1_0[22]_net_1\, 
        D => N_247, Y => \d_HADDR[22]\);
    
    \d_HADDR_0_iv[1]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \un13_d_haddr_1_m[1]\, B => 
        un46_d_haddr_cry_1_S, C => \d_HADDR_0_iv_1_0[1]_net_1\, D
         => N_247, Y => \d_HADDR[1]\);
    
    \HADDR_int[16]\ : SLE
      port map(D => \d_HADDR_0_iv_i_0[16]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[16]\);
    
    \state[9]\ : SLE
      port map(D => \state[10]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        HREADY_i_3_i_0, ALn => HPMS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[9]_net_1\);
    
    un13_d_haddr_1_cry_17 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[19]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_16\, S => un13_d_haddr_1_cry_17_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_17\);
    
    \d_ins2[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(13), B => un28_opcode, 
        Y => \d_ins2[13]_net_1\);
    
    \count_RNI2MQ7O[1]\ : CFG4
      generic map(INIT => x"EEAE")

      port map(A => \d_count_0_o3_3_0[1]\, B => 
        \d_count_0_a3_13_0[1]\, C => d_m2_e_1, D => 
        defSlaveSMNextState_m_0_3, Y => \d_count_0_o3_3_1[1]\);
    
    \bytecount[13]\ : SLE
      port map(D => N_52_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \bytecount[13]_net_1\);
    
    \haddr_write[13]\ : SLE
      port map(D => un46_d_haddr_cry_13_S, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_HWRITE_0_sqmuxa_1_0\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_write[13]_net_1\);
    
    state_21_rep1 : SLE
      port map(D => \state_ns_rep1[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state_21_rep1\);
    
    \rdata[28]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(28), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_725_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdata[28]_net_1\);
    
    \haddr_fetch[14]\ : SLE
      port map(D => N_2651_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_d_haddr_fetch_2_sqmuxa\, ALn => HPMS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \haddr_fetch[14]_net_1\);
    
    un1_state_44_0_12 : CFG4
      generic map(INIT => x"FEEE")

      port map(A => \un1_state_44_0_10\, B => N_4855, C => 
        HREADY_i_3, D => N_4827, Y => \un1_state_44_0_12\);
    
    un13_d_haddr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[10]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_7\, S => un13_d_haddr_1_cry_8_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_8\);
    
    \HWDATA_int[21]\ : SLE
      port map(D => \HWDATA_int_RNO[21]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(21));
    
    \haddr_fetch_RNO[23]\ : CFG4
      generic map(INIT => x"AAB8")

      port map(A => un13_d_haddr_1_cry_21_S, B => N_198, C => 
        \ConfigMaster_0_M_HADDR[23]\, D => N_4812, Y => 
        N_3216_i_0);
    
    \pause_count_RNO[2]\ : CFG3
      generic map(INIT => x"13")

      port map(A => N_66_i, B => N_3400, C => N_4813, Y => 
        N_4807_i_0);
    
    un46_d_haddr_cry_30 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[30]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un46_d_haddr_cry_29\, S => un46_d_haddr_cry_30_S, Y => 
        OPEN, FCO => \un46_d_haddr_cry_30\);
    
    \state_RNIADRJ[17]\ : CFG3
      generic map(INIT => x"0E")

      port map(A => \state[17]_net_1\, B => N_259, C => 
        HREADY_i_3, Y => N_725_i_0);
    
    d_HSIZE_1_sqmuxa_1_i_i_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => N_249, B => \state[24]_net_1\, Y => N_415);
    
    un1_state_46 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_state_42_0_0\, B => \un1_state_46_3\, Y
         => \un1_state_46\);
    
    \ins2[29]\ : SLE
      port map(D => \d_ins2[29]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[29]_net_1\);
    
    \expected[11]\ : SLE
      port map(D => ConfigMaster_0_M_HRDATA(11), CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_702_i_0, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \expected[11]_net_1\);
    
    \acc[7]\ : SLE
      port map(D => \d_acc[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \un1_state_25_0_0\, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \acc[7]_net_1\);
    
    \d_ins2[27]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ConfigMaster_0_M_HRDATA(27), B => un28_opcode, 
        Y => \d_ins2[27]_net_1\);
    
    \HADDR_int[5]\ : SLE
      port map(D => \d_HADDR[5]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_44_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ConfigMaster_0_M_HADDR[5]\);
    
    \state[26]\ : SLE
      port map(D => \state_ns[2]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \state[26]_net_1\);
    
    un13_d_haddr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \ConfigMaster_0_M_HADDR[4]\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un13_d_haddr_1_cry_1\, S => un13_d_haddr_1_cry_2_S, Y
         => OPEN, FCO => \un13_d_haddr_1_cry_2\);
    
    \d_HADDR_0_iv[23]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un1_d_HWRITE_0_sqmuxa_2, B => 
        \d_HADDR_0_iv_2[23]_net_1\, C => \haddr_fetch[23]_net_1\, 
        Y => \d_HADDR[23]\);
    
    \bytecount_RNO[5]\ : CFG3
      generic map(INIT => x"70")

      port map(A => \state[21]_net_1\, B => N_109_i, C => N_106, 
        Y => N_36_i_0);
    
    \ins2[17]\ : SLE
      port map(D => \d_ins2[17]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => N_654, ALn
         => HPMS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ins2[17]_net_1\);
    
    \HWDATA_int[20]\ : SLE
      port map(D => \HWDATA_int_RNO[20]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        un1_state_38_i_0, ALn => HPMS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => ConfigMaster_0_M_HWDATA(20));
    
    \d_acc[29]\ : CFG4
      generic map(INIT => x"EEE4")

      port map(A => \state[7]_net_1\, B => N_1166, C => 
        \ins2[29]_net_1\, D => \acc[29]_net_1\, Y => 
        \d_acc[29]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Igloo2_TFT_Video_Out_Test is

    port( MDDR_DQS                                : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                 : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DM_RDQS                            : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_BA                                 : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                               : out   std_logic_vector(15 downto 0);
          DEVRST_N                                : in    std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : out   std_logic;
          MDDR_WE_N                               : out   std_logic;
          MDDR_RESET_N                            : out   std_logic;
          MDDR_RAS_N                              : out   std_logic;
          MDDR_ODT                                : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                   : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                    : in    std_logic;
          MDDR_CS_N                               : out   std_logic;
          MDDR_CKE                                : out   std_logic;
          MDDR_CAS_N                              : out   std_logic;
          MDDR_CLK_N                              : out   std_logic;
          MDDR_CLK                                : out   std_logic
        );

end Igloo2_TFT_Video_Out_Test;

architecture DEF_ARCH of Igloo2_TFT_Video_Out_Test is 

  component Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_O2F                        : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreResetP
    port( HPMS_READY                                       : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F                      : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0          : in    std_logic := 'U';
          INIT_DONE                                        : out   std_logic;
          POWER_ON_RESET_N                                 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic := 'U';
          CORECONFIGP_0_CONFIG1_DONE                       : in    std_logic := 'U';
          CORECONFIGP_0_CONFIG2_DONE                       : in    std_logic := 'U';
          CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET     : in    std_logic := 'U';
          CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N         : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component Igloo2_TFT_Video_Out_Test_HPMS
    port( MDDR_DQS                                                    : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                                     : inout   std_logic_vector(15 downto 0);
          MDDR_DM_RDQS                                                : inout   std_logic_vector(1 downto 0);
          MDDR_BA                                                     : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                                   : out   std_logic_vector(15 downto 0);
          xhdl1328_i_m_0_1                                            : in    std_logic_vector(0 to 0) := (others => 'U');
          ConfigMaster_0_M_HRDATA                                     : out   std_logic_vector(31 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA                         : out   std_logic_vector(15 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HSIZE                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HTRANS                            : in    std_logic_vector(1 to 1) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HWDATA                            : in    std_logic_vector(31 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR                          : in    std_logic_vector(10 downto 2) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PWDATA                         : in    std_logic_vector(15 downto 0) := (others => 'U');
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_0  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_1  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_2  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_3  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_4  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_5  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_6  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_7  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_8  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_9  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_10 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_11 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_12 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_13 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_14 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_15 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_16 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18 : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N                                : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                                    : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i_0                                : out   std_logic;
          MDDR_WE_N                                                   : out   std_logic;
          MDDR_RESET_N                                                : out   std_logic;
          MDDR_RAS_N                                                  : out   std_logic;
          MDDR_ODT                                                    : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                                       : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                                        : in    std_logic := 'U';
          MDDR_CS_N                                                   : out   std_logic;
          MDDR_CKE                                                    : out   std_logic;
          MDDR_CAS_N                                                  : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY                            : inout   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m                        : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F            : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE   : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx     : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE    : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY                         : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR                        : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HSELx                             : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HWRITE                            : in    std_logic := 'U';
          HPMS_DDR_FIC_SUBSYSTEM_LOCK                                 : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY    : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR   : in    std_logic := 'U';
          CORECONFIGP_0_SOFT_RESET_F2M_i_0                            : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0                     : in    std_logic := 'U';
          CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N                    : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE                        : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx                          : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PWRITE                         : in    std_logic := 'U';
          MDDR_CLK_N                                                  : out   std_logic;
          MDDR_CLK                                                    : out   std_logic
        );
  end component;

  component Igloo2_TFT_Video_Out_Test_CCC_0_FCCC
    port( Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0            : out   std_logic;
          HPMS_DDR_FIC_SUBSYSTEM_LOCK                        : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CoreConfigP
    port( Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA    : in    std_logic_vector(16 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PWDATA                         : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR                          : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA                         : in    std_logic_vector(15 downto 0) := (others => 'U');
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9  : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18 : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11  : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13  : in    std_logic := 'U';
          CORECONFIGP_0_SOFT_RESET_F2M_i_0                            : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY    : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                                : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PCLK                                    : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR   : out   std_logic;
          CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET                : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                                  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                                  : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE                         : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE    : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PCLK_i_0                                : in    std_logic := 'U';
          INIT_DONE                                                   : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE                        : out   std_logic;
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE   : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx     : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx                          : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR                        : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PREADY                         : in    std_logic := 'U'
        );
  end component;

  component 
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0
    port( ConfigMaster_0_M_HSIZE                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          ConfigMaster_0_M_HADDR                  : in    std_logic_vector(31 downto 0) := (others => 'U');
          ConfigMaster_0_M_HTRANS                 : in    std_logic_vector(1 to 1) := (others => 'U');
          xhdl1328_i_m_0_1                        : out   std_logic_vector(0 to 0);
          masterDataInProg                        : out   std_logic_vector(0 to 0);
          ConfigMaster_0_M_HWDATA                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_1_AHBmslave16_HWDATA        : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HSIZE         : out   std_logic_vector(1 downto 0);
          CoreAHBLite_1_AHBmslave16_HADDR         : out   std_logic_vector(31 downto 0);
          CoreAHBLite_1_AHBmslave16_HTRANS        : out   std_logic_vector(1 to 1);
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          ConfigMaster_0_M_HWRITE                 : in    std_logic := 'U';
          defSlaveSMNextState_m_0_3               : out   std_logic;
          un1_state_31_i_i_a2_0_d_1_0_1           : out   std_logic;
          defSlaveSMNextState_m_0_2               : out   std_logic;
          HREADY_i_3                              : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : out   std_logic;
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : out   std_logic;
          N_98                                    : out   std_logic;
          N_25                                    : out   std_logic;
          defSlaveSMNextState_m_0_3_1             : out   std_logic;
          defSlaveSMNextState_m                   : out   std_logic;
          HREADY_i_3_i_0                          : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HREADY_i_m    : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HSELx         : out   std_logic;
          CoreAHBLite_1_AHBmslave16_HWRITE        : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component CoreConfigMaster
    port( ConfigMaster_0_M_HTRANS                 : out   std_logic_vector(1 to 1);
          ConfigMaster_0_M_HWDATA                 : out   std_logic_vector(31 downto 0);
          ConfigMaster_0_M_HSIZE                  : out   std_logic_vector(1 downto 0);
          ConfigMaster_0_M_HRDATA                 : in    std_logic_vector(31 downto 0) := (others => 'U');
          ConfigMaster_0_M_HADDR                  : out   std_logic_vector(31 downto 0);
          masterDataInProg                        : in    std_logic_vector(0 to 0) := (others => 'U');
          xhdl1328_i_m_0_1                        : in    std_logic_vector(0 to 0) := (others => 'U');
          HPMS_READY                              : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          ConfigMaster_0_M_HWRITE                 : out   std_logic;
          HREADY_i_3_i_0                          : in    std_logic := 'U';
          defSlaveSMNextState_m_0_3               : in    std_logic := 'U';
          defSlaveSMNextState_m_0_2               : in    std_logic := 'U';
          CoreAHBLite_1_AHBmslave16_HREADY        : in    std_logic := 'U';
          defSlaveSMNextState_m                   : in    std_logic := 'U';
          HREADY_i_3                              : in    std_logic := 'U';
          un1_state_31_i_i_a2_0_d_1_0_1           : in    std_logic := 'U';
          defSlaveSMNextState_i_a2_0_RNI3J724_2   : in    std_logic := 'U';
          defSlaveSMNextState_i_a2_0_RNI3J724_1   : in    std_logic := 'U';
          N_98                                    : in    std_logic := 'U';
          N_25                                    : in    std_logic := 'U';
          defSlaveSMNextState_m_0_3_1             : in    std_logic := 'U'
        );
  end component;

    signal POWER_ON_RESET_N, 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \ConfigMaster_0_M_HTRANS[1]\, 
        \ConfigMaster_0_M_HWDATA[0]\, 
        \ConfigMaster_0_M_HWDATA[1]\, 
        \ConfigMaster_0_M_HWDATA[2]\, 
        \ConfigMaster_0_M_HWDATA[3]\, 
        \ConfigMaster_0_M_HWDATA[4]\, 
        \ConfigMaster_0_M_HWDATA[5]\, 
        \ConfigMaster_0_M_HWDATA[6]\, 
        \ConfigMaster_0_M_HWDATA[7]\, 
        \ConfigMaster_0_M_HWDATA[8]\, 
        \ConfigMaster_0_M_HWDATA[9]\, 
        \ConfigMaster_0_M_HWDATA[10]\, 
        \ConfigMaster_0_M_HWDATA[11]\, 
        \ConfigMaster_0_M_HWDATA[12]\, 
        \ConfigMaster_0_M_HWDATA[13]\, 
        \ConfigMaster_0_M_HWDATA[14]\, 
        \ConfigMaster_0_M_HWDATA[15]\, 
        \ConfigMaster_0_M_HWDATA[16]\, 
        \ConfigMaster_0_M_HWDATA[17]\, 
        \ConfigMaster_0_M_HWDATA[18]\, 
        \ConfigMaster_0_M_HWDATA[19]\, 
        \ConfigMaster_0_M_HWDATA[20]\, 
        \ConfigMaster_0_M_HWDATA[21]\, 
        \ConfigMaster_0_M_HWDATA[22]\, 
        \ConfigMaster_0_M_HWDATA[23]\, 
        \ConfigMaster_0_M_HWDATA[24]\, 
        \ConfigMaster_0_M_HWDATA[25]\, 
        \ConfigMaster_0_M_HWDATA[26]\, 
        \ConfigMaster_0_M_HWDATA[27]\, 
        \ConfigMaster_0_M_HWDATA[28]\, 
        \ConfigMaster_0_M_HWDATA[29]\, 
        \ConfigMaster_0_M_HWDATA[30]\, 
        \ConfigMaster_0_M_HWDATA[31]\, 
        \ConfigMaster_0_M_HSIZE[0]\, \ConfigMaster_0_M_HSIZE[1]\, 
        \ConfigMaster_0_M_HRDATA[0]\, 
        \ConfigMaster_0_M_HRDATA[1]\, 
        \ConfigMaster_0_M_HRDATA[2]\, 
        \ConfigMaster_0_M_HRDATA[3]\, 
        \ConfigMaster_0_M_HRDATA[4]\, 
        \ConfigMaster_0_M_HRDATA[5]\, 
        \ConfigMaster_0_M_HRDATA[6]\, 
        \ConfigMaster_0_M_HRDATA[7]\, 
        \ConfigMaster_0_M_HRDATA[8]\, 
        \ConfigMaster_0_M_HRDATA[9]\, 
        \ConfigMaster_0_M_HRDATA[10]\, 
        \ConfigMaster_0_M_HRDATA[11]\, 
        \ConfigMaster_0_M_HRDATA[12]\, 
        \ConfigMaster_0_M_HRDATA[13]\, 
        \ConfigMaster_0_M_HRDATA[14]\, 
        \ConfigMaster_0_M_HRDATA[15]\, 
        \ConfigMaster_0_M_HRDATA[16]\, 
        \ConfigMaster_0_M_HRDATA[17]\, 
        \ConfigMaster_0_M_HRDATA[18]\, 
        \ConfigMaster_0_M_HRDATA[19]\, 
        \ConfigMaster_0_M_HRDATA[20]\, 
        \ConfigMaster_0_M_HRDATA[21]\, 
        \ConfigMaster_0_M_HRDATA[22]\, 
        \ConfigMaster_0_M_HRDATA[23]\, 
        \ConfigMaster_0_M_HRDATA[24]\, 
        \ConfigMaster_0_M_HRDATA[25]\, 
        \ConfigMaster_0_M_HRDATA[26]\, 
        \ConfigMaster_0_M_HRDATA[27]\, 
        \ConfigMaster_0_M_HRDATA[28]\, 
        \ConfigMaster_0_M_HRDATA[29]\, 
        \ConfigMaster_0_M_HRDATA[30]\, 
        \ConfigMaster_0_M_HRDATA[31]\, 
        \ConfigMaster_0_M_HADDR[0]\, \ConfigMaster_0_M_HADDR[1]\, 
        \ConfigMaster_0_M_HADDR[2]\, \ConfigMaster_0_M_HADDR[3]\, 
        \ConfigMaster_0_M_HADDR[4]\, \ConfigMaster_0_M_HADDR[5]\, 
        \ConfigMaster_0_M_HADDR[6]\, \ConfigMaster_0_M_HADDR[7]\, 
        \ConfigMaster_0_M_HADDR[8]\, \ConfigMaster_0_M_HADDR[9]\, 
        \ConfigMaster_0_M_HADDR[10]\, 
        \ConfigMaster_0_M_HADDR[11]\, 
        \ConfigMaster_0_M_HADDR[12]\, 
        \ConfigMaster_0_M_HADDR[13]\, 
        \ConfigMaster_0_M_HADDR[14]\, 
        \ConfigMaster_0_M_HADDR[15]\, 
        \ConfigMaster_0_M_HADDR[16]\, 
        \ConfigMaster_0_M_HADDR[17]\, 
        \ConfigMaster_0_M_HADDR[18]\, 
        \ConfigMaster_0_M_HADDR[19]\, 
        \ConfigMaster_0_M_HADDR[20]\, 
        \ConfigMaster_0_M_HADDR[21]\, 
        \ConfigMaster_0_M_HADDR[22]\, 
        \ConfigMaster_0_M_HADDR[23]\, 
        \ConfigMaster_0_M_HADDR[24]\, 
        \ConfigMaster_0_M_HADDR[25]\, 
        \ConfigMaster_0_M_HADDR[26]\, 
        \ConfigMaster_0_M_HADDR[27]\, 
        \ConfigMaster_0_M_HADDR[28]\, 
        \ConfigMaster_0_M_HADDR[29]\, 
        \ConfigMaster_0_M_HADDR[30]\, 
        \ConfigMaster_0_M_HADDR[31]\, \masterDataInProg[0]\, 
        \xhdl1328_i_m_0_1[0]\, HPMS_READY, 
        ConfigMaster_0_M_HWRITE, HREADY_i_3_i_0, 
        defSlaveSMNextState_m_0_3, defSlaveSMNextState_m_0_2, 
        CoreAHBLite_1_AHBmslave16_HREADY, defSlaveSMNextState_m, 
        HREADY_i_3, un1_state_31_i_i_a2_0_d_1_0_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, N_98, N_25, 
        defSlaveSMNextState_m_0_3_1, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[0]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[1]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[2]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[3]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[4]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[5]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[6]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[7]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[8]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[9]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[10]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[11]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[12]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[13]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[14]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[15]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[16]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[17]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[18]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[19]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[20]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[21]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[22]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[23]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[24]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[25]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[26]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[27]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[28]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[29]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[30]\, 
        \CoreAHBLite_1_AHBmslave16_HWDATA[31]\, 
        \CoreAHBLite_1_AHBmslave16_HSIZE[0]\, 
        \CoreAHBLite_1_AHBmslave16_HSIZE[1]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[0]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[1]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[2]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[3]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[4]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[5]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[6]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[7]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[8]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[9]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[10]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[11]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[12]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[13]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[14]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[15]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[16]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[17]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[18]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[19]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[20]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[21]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[22]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[23]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[24]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[25]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[26]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[27]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[28]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[29]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[30]\, 
        \CoreAHBLite_1_AHBmslave16_HADDR[31]\, 
        \CoreAHBLite_1_AHBmslave16_HTRANS[1]\, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, 
        CoreAHBLite_1_AHBmslave16_HSELx, 
        CoreAHBLite_1_AHBmslave16_HWRITE, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[18]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[2]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[3]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[4]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[5]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[6]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[7]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[8]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[9]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[10]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[12]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[13]\, 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[15]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_APB_S_PRESET_N, CORECONFIGP_0_APB_S_PCLK, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR, 
        CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET, 
        CORECONFIGP_0_CONFIG1_DONE, CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_APB_S_PCLK_i_0, INIT_DONE, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        FABOSC_0_RCOSC_25_50MHZ_O2F, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N, GND_net_1, 
        VCC_net_1 : std_logic;

    for all : Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC
	Use entity work.Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : Igloo2_TFT_Video_Out_Test_HPMS
	Use entity work.Igloo2_TFT_Video_Out_Test_HPMS(DEF_ARCH);
    for all : Igloo2_TFT_Video_Out_Test_CCC_0_FCCC
	Use entity work.Igloo2_TFT_Video_Out_Test_CCC_0_FCCC(DEF_ARCH);
    for all : CoreConfigP
	Use entity work.CoreConfigP(DEF_ARCH);
    for all : CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0
	Use entity work.
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0(DEF_ARCH);
    for all : CoreConfigMaster
	Use entity work.CoreConfigMaster(DEF_ARCH);
begin 

    Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 <= 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\;

    FABOSC_0 : Igloo2_TFT_Video_Out_Test_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CORERESETP_0 : CoreResetP
      port map(HPMS_READY => HPMS_READY, 
        FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, INIT_DONE => 
        INIT_DONE, POWER_ON_RESET_N => POWER_ON_RESET_N, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, CORECONFIGP_0_CONFIG1_DONE
         => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_CONFIG2_DONE => CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET => 
        CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET, 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N => 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    Igloo2_TFT_Video_Out_Test_HPMS_0 : 
        Igloo2_TFT_Video_Out_Test_HPMS
      port map(MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14) => 
        MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12) => 
        MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10) => 
        MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), 
        MDDR_DM_RDQS(0) => MDDR_DM_RDQS(0), MDDR_BA(2) => 
        MDDR_BA(2), MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => 
        MDDR_BA(0), MDDR_ADDR(15) => MDDR_ADDR(15), MDDR_ADDR(14)
         => MDDR_ADDR(14), MDDR_ADDR(13) => MDDR_ADDR(13), 
        MDDR_ADDR(12) => MDDR_ADDR(12), MDDR_ADDR(11) => 
        MDDR_ADDR(11), MDDR_ADDR(10) => MDDR_ADDR(10), 
        MDDR_ADDR(9) => MDDR_ADDR(9), MDDR_ADDR(8) => 
        MDDR_ADDR(8), MDDR_ADDR(7) => MDDR_ADDR(7), MDDR_ADDR(6)
         => MDDR_ADDR(6), MDDR_ADDR(5) => MDDR_ADDR(5), 
        MDDR_ADDR(4) => MDDR_ADDR(4), MDDR_ADDR(3) => 
        MDDR_ADDR(3), MDDR_ADDR(2) => MDDR_ADDR(2), MDDR_ADDR(1)
         => MDDR_ADDR(1), MDDR_ADDR(0) => MDDR_ADDR(0), 
        xhdl1328_i_m_0_1(0) => \xhdl1328_i_m_0_1[0]\, 
        ConfigMaster_0_M_HRDATA(31) => 
        \ConfigMaster_0_M_HRDATA[31]\, 
        ConfigMaster_0_M_HRDATA(30) => 
        \ConfigMaster_0_M_HRDATA[30]\, 
        ConfigMaster_0_M_HRDATA(29) => 
        \ConfigMaster_0_M_HRDATA[29]\, 
        ConfigMaster_0_M_HRDATA(28) => 
        \ConfigMaster_0_M_HRDATA[28]\, 
        ConfigMaster_0_M_HRDATA(27) => 
        \ConfigMaster_0_M_HRDATA[27]\, 
        ConfigMaster_0_M_HRDATA(26) => 
        \ConfigMaster_0_M_HRDATA[26]\, 
        ConfigMaster_0_M_HRDATA(25) => 
        \ConfigMaster_0_M_HRDATA[25]\, 
        ConfigMaster_0_M_HRDATA(24) => 
        \ConfigMaster_0_M_HRDATA[24]\, 
        ConfigMaster_0_M_HRDATA(23) => 
        \ConfigMaster_0_M_HRDATA[23]\, 
        ConfigMaster_0_M_HRDATA(22) => 
        \ConfigMaster_0_M_HRDATA[22]\, 
        ConfigMaster_0_M_HRDATA(21) => 
        \ConfigMaster_0_M_HRDATA[21]\, 
        ConfigMaster_0_M_HRDATA(20) => 
        \ConfigMaster_0_M_HRDATA[20]\, 
        ConfigMaster_0_M_HRDATA(19) => 
        \ConfigMaster_0_M_HRDATA[19]\, 
        ConfigMaster_0_M_HRDATA(18) => 
        \ConfigMaster_0_M_HRDATA[18]\, 
        ConfigMaster_0_M_HRDATA(17) => 
        \ConfigMaster_0_M_HRDATA[17]\, 
        ConfigMaster_0_M_HRDATA(16) => 
        \ConfigMaster_0_M_HRDATA[16]\, 
        ConfigMaster_0_M_HRDATA(15) => 
        \ConfigMaster_0_M_HRDATA[15]\, 
        ConfigMaster_0_M_HRDATA(14) => 
        \ConfigMaster_0_M_HRDATA[14]\, 
        ConfigMaster_0_M_HRDATA(13) => 
        \ConfigMaster_0_M_HRDATA[13]\, 
        ConfigMaster_0_M_HRDATA(12) => 
        \ConfigMaster_0_M_HRDATA[12]\, 
        ConfigMaster_0_M_HRDATA(11) => 
        \ConfigMaster_0_M_HRDATA[11]\, 
        ConfigMaster_0_M_HRDATA(10) => 
        \ConfigMaster_0_M_HRDATA[10]\, ConfigMaster_0_M_HRDATA(9)
         => \ConfigMaster_0_M_HRDATA[9]\, 
        ConfigMaster_0_M_HRDATA(8) => 
        \ConfigMaster_0_M_HRDATA[8]\, ConfigMaster_0_M_HRDATA(7)
         => \ConfigMaster_0_M_HRDATA[7]\, 
        ConfigMaster_0_M_HRDATA(6) => 
        \ConfigMaster_0_M_HRDATA[6]\, ConfigMaster_0_M_HRDATA(5)
         => \ConfigMaster_0_M_HRDATA[5]\, 
        ConfigMaster_0_M_HRDATA(4) => 
        \ConfigMaster_0_M_HRDATA[4]\, ConfigMaster_0_M_HRDATA(3)
         => \ConfigMaster_0_M_HRDATA[3]\, 
        ConfigMaster_0_M_HRDATA(2) => 
        \ConfigMaster_0_M_HRDATA[2]\, ConfigMaster_0_M_HRDATA(1)
         => \ConfigMaster_0_M_HRDATA[1]\, 
        ConfigMaster_0_M_HRDATA(0) => 
        \ConfigMaster_0_M_HRDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(31) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[31]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(30) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[30]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(29) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[29]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(28) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[28]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(27) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[27]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(26) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[26]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(25) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[25]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(24) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[24]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(23) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[23]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(22) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[22]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(21) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[21]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(20) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[20]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(19) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[19]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(18) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[18]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(17) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[17]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(16) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[16]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(15) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[15]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(14) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[14]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(13) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[13]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(12) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[12]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(11) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[11]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(10) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[10]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(9) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[9]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(8) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[8]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(7) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[7]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(6) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[6]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(5) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[5]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(4) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[4]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(3) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[3]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(2) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[2]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(1) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[1]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(0) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[0]\, 
        CoreAHBLite_1_AHBmslave16_HSIZE(1) => 
        \CoreAHBLite_1_AHBmslave16_HSIZE[1]\, 
        CoreAHBLite_1_AHBmslave16_HSIZE(0) => 
        \CoreAHBLite_1_AHBmslave16_HSIZE[0]\, 
        CoreAHBLite_1_AHBmslave16_HTRANS(1) => 
        \CoreAHBLite_1_AHBmslave16_HTRANS[1]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(31) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[31]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(30) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[30]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(29) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[29]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(28) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[28]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(27) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[27]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(26) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[26]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(25) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[25]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(24) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[24]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(23) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[23]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(22) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[22]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(21) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[21]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(20) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[20]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(19) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[19]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(18) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[18]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(17) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[17]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(16) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[16]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(15) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[15]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(14) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[14]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(13) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[13]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(12) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[12]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(11) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[11]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(10) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[10]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(9) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[9]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(8) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[8]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(7) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[7]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(6) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[6]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(5) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[5]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(4) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[4]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(3) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[3]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(2) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[2]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(1) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[1]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(0) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[15]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_0
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_1
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_2
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_3
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_4
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_5
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_6
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_7
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_8
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_9
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_10
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_11
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_12
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_13
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_14
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_15
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA_16
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[18]\, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, CORECONFIGP_0_APB_S_PCLK
         => CORECONFIGP_0_APB_S_PCLK, 
        CORECONFIGP_0_APB_S_PCLK_i_0 => 
        CORECONFIGP_0_APB_S_PCLK_i_0, MDDR_WE_N => MDDR_WE_N, 
        MDDR_RESET_N => MDDR_RESET_N, MDDR_RAS_N => MDDR_RAS_N, 
        MDDR_ODT => MDDR_ODT, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_CS_N => MDDR_CS_N, MDDR_CKE
         => MDDR_CKE, MDDR_CAS_N => MDDR_CAS_N, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_MSS_RESET_N_M2F, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CoreAHBLite_1_AHBmslave16_HSELx => 
        CoreAHBLite_1_AHBmslave16_HSELx, 
        CoreAHBLite_1_AHBmslave16_HWRITE => 
        CoreAHBLite_1_AHBmslave16_HWRITE, 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK => 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR, 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0 => 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N => 
        CORERESETP_0_MDDR_DDR_AXI_S_CORE_RESET_N, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, MDDR_CLK_N => 
        MDDR_CLK_N, MDDR_CLK => MDDR_CLK);
    
    CCC_0 : Igloo2_TFT_Video_Out_Test_CCC_0_FCCC
      port map(Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK => 
        HPMS_DDR_FIC_SUBSYSTEM_LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CORECONFIGP_0 : CoreConfigP
      port map(
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(16)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(15)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(14)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(13)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(12)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(11)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(10)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(9)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(8)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(7)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(6)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(5)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(4)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(3)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(2)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(1)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA(0)
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_0
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_1
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_2
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_3
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_4
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_5
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_6
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_7
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_8
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_9
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_10
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_11
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_12
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_13
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_14
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_15
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_16
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA_18
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PRDATA[18]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_0
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[2]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_1
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[3]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_2
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[4]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_3
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[5]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_4
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[6]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_5
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[7]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_6
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[8]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_7
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[9]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_8
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[10]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_10
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[12]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_11
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[13]\, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR_13
         => 
        \Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PADDR[15]\, 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0 => 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, CORECONFIGP_0_APB_S_PCLK
         => CORECONFIGP_0_APB_S_PCLK, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSLVERR, 
        CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET => 
        CORECONFIGP_0_SOFT_MDDR_DDR_AXI_S_CORE_RESET, 
        CORECONFIGP_0_CONFIG1_DONE => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_CONFIG2_DONE => CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_APB_S_PCLK_i_0 => 
        CORECONFIGP_0_APB_S_PCLK_i_0, INIT_DONE => INIT_DONE, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PENABLE, 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx
         => 
        Igloo2_TFT_Video_Out_Test_HPMS_0_FIC_2_APB_MASTER_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY);
    
    CoreAHBLite_1 : 
        CoreAHBLite_19_1_1_1_0_1_0_1_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0
      port map(ConfigMaster_0_M_HSIZE(1) => 
        \ConfigMaster_0_M_HSIZE[1]\, ConfigMaster_0_M_HSIZE(0)
         => \ConfigMaster_0_M_HSIZE[0]\, 
        ConfigMaster_0_M_HADDR(31) => 
        \ConfigMaster_0_M_HADDR[31]\, ConfigMaster_0_M_HADDR(30)
         => \ConfigMaster_0_M_HADDR[30]\, 
        ConfigMaster_0_M_HADDR(29) => 
        \ConfigMaster_0_M_HADDR[29]\, ConfigMaster_0_M_HADDR(28)
         => \ConfigMaster_0_M_HADDR[28]\, 
        ConfigMaster_0_M_HADDR(27) => 
        \ConfigMaster_0_M_HADDR[27]\, ConfigMaster_0_M_HADDR(26)
         => \ConfigMaster_0_M_HADDR[26]\, 
        ConfigMaster_0_M_HADDR(25) => 
        \ConfigMaster_0_M_HADDR[25]\, ConfigMaster_0_M_HADDR(24)
         => \ConfigMaster_0_M_HADDR[24]\, 
        ConfigMaster_0_M_HADDR(23) => 
        \ConfigMaster_0_M_HADDR[23]\, ConfigMaster_0_M_HADDR(22)
         => \ConfigMaster_0_M_HADDR[22]\, 
        ConfigMaster_0_M_HADDR(21) => 
        \ConfigMaster_0_M_HADDR[21]\, ConfigMaster_0_M_HADDR(20)
         => \ConfigMaster_0_M_HADDR[20]\, 
        ConfigMaster_0_M_HADDR(19) => 
        \ConfigMaster_0_M_HADDR[19]\, ConfigMaster_0_M_HADDR(18)
         => \ConfigMaster_0_M_HADDR[18]\, 
        ConfigMaster_0_M_HADDR(17) => 
        \ConfigMaster_0_M_HADDR[17]\, ConfigMaster_0_M_HADDR(16)
         => \ConfigMaster_0_M_HADDR[16]\, 
        ConfigMaster_0_M_HADDR(15) => 
        \ConfigMaster_0_M_HADDR[15]\, ConfigMaster_0_M_HADDR(14)
         => \ConfigMaster_0_M_HADDR[14]\, 
        ConfigMaster_0_M_HADDR(13) => 
        \ConfigMaster_0_M_HADDR[13]\, ConfigMaster_0_M_HADDR(12)
         => \ConfigMaster_0_M_HADDR[12]\, 
        ConfigMaster_0_M_HADDR(11) => 
        \ConfigMaster_0_M_HADDR[11]\, ConfigMaster_0_M_HADDR(10)
         => \ConfigMaster_0_M_HADDR[10]\, 
        ConfigMaster_0_M_HADDR(9) => \ConfigMaster_0_M_HADDR[9]\, 
        ConfigMaster_0_M_HADDR(8) => \ConfigMaster_0_M_HADDR[8]\, 
        ConfigMaster_0_M_HADDR(7) => \ConfigMaster_0_M_HADDR[7]\, 
        ConfigMaster_0_M_HADDR(6) => \ConfigMaster_0_M_HADDR[6]\, 
        ConfigMaster_0_M_HADDR(5) => \ConfigMaster_0_M_HADDR[5]\, 
        ConfigMaster_0_M_HADDR(4) => \ConfigMaster_0_M_HADDR[4]\, 
        ConfigMaster_0_M_HADDR(3) => \ConfigMaster_0_M_HADDR[3]\, 
        ConfigMaster_0_M_HADDR(2) => \ConfigMaster_0_M_HADDR[2]\, 
        ConfigMaster_0_M_HADDR(1) => \ConfigMaster_0_M_HADDR[1]\, 
        ConfigMaster_0_M_HADDR(0) => \ConfigMaster_0_M_HADDR[0]\, 
        ConfigMaster_0_M_HTRANS(1) => 
        \ConfigMaster_0_M_HTRANS[1]\, xhdl1328_i_m_0_1(0) => 
        \xhdl1328_i_m_0_1[0]\, masterDataInProg(0) => 
        \masterDataInProg[0]\, ConfigMaster_0_M_HWDATA(31) => 
        \ConfigMaster_0_M_HWDATA[31]\, 
        ConfigMaster_0_M_HWDATA(30) => 
        \ConfigMaster_0_M_HWDATA[30]\, 
        ConfigMaster_0_M_HWDATA(29) => 
        \ConfigMaster_0_M_HWDATA[29]\, 
        ConfigMaster_0_M_HWDATA(28) => 
        \ConfigMaster_0_M_HWDATA[28]\, 
        ConfigMaster_0_M_HWDATA(27) => 
        \ConfigMaster_0_M_HWDATA[27]\, 
        ConfigMaster_0_M_HWDATA(26) => 
        \ConfigMaster_0_M_HWDATA[26]\, 
        ConfigMaster_0_M_HWDATA(25) => 
        \ConfigMaster_0_M_HWDATA[25]\, 
        ConfigMaster_0_M_HWDATA(24) => 
        \ConfigMaster_0_M_HWDATA[24]\, 
        ConfigMaster_0_M_HWDATA(23) => 
        \ConfigMaster_0_M_HWDATA[23]\, 
        ConfigMaster_0_M_HWDATA(22) => 
        \ConfigMaster_0_M_HWDATA[22]\, 
        ConfigMaster_0_M_HWDATA(21) => 
        \ConfigMaster_0_M_HWDATA[21]\, 
        ConfigMaster_0_M_HWDATA(20) => 
        \ConfigMaster_0_M_HWDATA[20]\, 
        ConfigMaster_0_M_HWDATA(19) => 
        \ConfigMaster_0_M_HWDATA[19]\, 
        ConfigMaster_0_M_HWDATA(18) => 
        \ConfigMaster_0_M_HWDATA[18]\, 
        ConfigMaster_0_M_HWDATA(17) => 
        \ConfigMaster_0_M_HWDATA[17]\, 
        ConfigMaster_0_M_HWDATA(16) => 
        \ConfigMaster_0_M_HWDATA[16]\, 
        ConfigMaster_0_M_HWDATA(15) => 
        \ConfigMaster_0_M_HWDATA[15]\, 
        ConfigMaster_0_M_HWDATA(14) => 
        \ConfigMaster_0_M_HWDATA[14]\, 
        ConfigMaster_0_M_HWDATA(13) => 
        \ConfigMaster_0_M_HWDATA[13]\, 
        ConfigMaster_0_M_HWDATA(12) => 
        \ConfigMaster_0_M_HWDATA[12]\, 
        ConfigMaster_0_M_HWDATA(11) => 
        \ConfigMaster_0_M_HWDATA[11]\, 
        ConfigMaster_0_M_HWDATA(10) => 
        \ConfigMaster_0_M_HWDATA[10]\, ConfigMaster_0_M_HWDATA(9)
         => \ConfigMaster_0_M_HWDATA[9]\, 
        ConfigMaster_0_M_HWDATA(8) => 
        \ConfigMaster_0_M_HWDATA[8]\, ConfigMaster_0_M_HWDATA(7)
         => \ConfigMaster_0_M_HWDATA[7]\, 
        ConfigMaster_0_M_HWDATA(6) => 
        \ConfigMaster_0_M_HWDATA[6]\, ConfigMaster_0_M_HWDATA(5)
         => \ConfigMaster_0_M_HWDATA[5]\, 
        ConfigMaster_0_M_HWDATA(4) => 
        \ConfigMaster_0_M_HWDATA[4]\, ConfigMaster_0_M_HWDATA(3)
         => \ConfigMaster_0_M_HWDATA[3]\, 
        ConfigMaster_0_M_HWDATA(2) => 
        \ConfigMaster_0_M_HWDATA[2]\, ConfigMaster_0_M_HWDATA(1)
         => \ConfigMaster_0_M_HWDATA[1]\, 
        ConfigMaster_0_M_HWDATA(0) => 
        \ConfigMaster_0_M_HWDATA[0]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(31) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[31]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(30) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[30]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(29) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[29]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(28) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[28]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(27) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[27]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(26) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[26]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(25) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[25]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(24) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[24]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(23) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[23]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(22) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[22]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(21) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[21]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(20) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[20]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(19) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[19]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(18) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[18]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(17) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[17]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(16) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[16]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(15) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[15]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(14) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[14]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(13) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[13]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(12) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[12]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(11) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[11]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(10) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[10]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(9) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[9]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(8) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[8]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(7) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[7]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(6) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[6]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(5) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[5]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(4) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[4]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(3) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[3]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(2) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[2]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(1) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[1]\, 
        CoreAHBLite_1_AHBmslave16_HWDATA(0) => 
        \CoreAHBLite_1_AHBmslave16_HWDATA[0]\, 
        CoreAHBLite_1_AHBmslave16_HSIZE(1) => 
        \CoreAHBLite_1_AHBmslave16_HSIZE[1]\, 
        CoreAHBLite_1_AHBmslave16_HSIZE(0) => 
        \CoreAHBLite_1_AHBmslave16_HSIZE[0]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(31) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[31]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(30) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[30]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(29) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[29]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(28) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[28]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(27) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[27]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(26) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[26]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(25) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[25]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(24) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[24]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(23) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[23]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(22) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[22]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(21) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[21]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(20) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[20]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(19) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[19]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(18) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[18]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(17) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[17]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(16) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[16]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(15) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[15]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(14) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[14]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(13) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[13]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(12) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[12]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(11) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[11]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(10) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[10]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(9) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[9]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(8) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[8]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(7) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[7]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(6) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[6]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(5) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[5]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(4) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[4]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(3) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[3]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(2) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[2]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(1) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[1]\, 
        CoreAHBLite_1_AHBmslave16_HADDR(0) => 
        \CoreAHBLite_1_AHBmslave16_HADDR[0]\, 
        CoreAHBLite_1_AHBmslave16_HTRANS(1) => 
        \CoreAHBLite_1_AHBmslave16_HTRANS[1]\, HPMS_READY => 
        HPMS_READY, Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, 
        ConfigMaster_0_M_HWRITE => ConfigMaster_0_M_HWRITE, 
        defSlaveSMNextState_m_0_3 => defSlaveSMNextState_m_0_3, 
        un1_state_31_i_i_a2_0_d_1_0_1 => 
        un1_state_31_i_i_a2_0_d_1_0_1, defSlaveSMNextState_m_0_2
         => defSlaveSMNextState_m_0_2, HREADY_i_3 => HREADY_i_3, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, N_98 => N_98, N_25
         => N_25, defSlaveSMNextState_m_0_3_1 => 
        defSlaveSMNextState_m_0_3_1, defSlaveSMNextState_m => 
        defSlaveSMNextState_m, HREADY_i_3_i_0 => HREADY_i_3_i_0, 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m => 
        CoreAHBLite_1_AHBmslave16_HREADY_i_m, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, 
        CoreAHBLite_1_AHBmslave16_HSELx => 
        CoreAHBLite_1_AHBmslave16_HSELx, 
        CoreAHBLite_1_AHBmslave16_HWRITE => 
        CoreAHBLite_1_AHBmslave16_HWRITE);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => POWER_ON_RESET_N, DEVRST_N => 
        DEVRST_N);
    
    ConfigMaster_0 : CoreConfigMaster
      port map(ConfigMaster_0_M_HTRANS(1) => 
        \ConfigMaster_0_M_HTRANS[1]\, ConfigMaster_0_M_HWDATA(31)
         => \ConfigMaster_0_M_HWDATA[31]\, 
        ConfigMaster_0_M_HWDATA(30) => 
        \ConfigMaster_0_M_HWDATA[30]\, 
        ConfigMaster_0_M_HWDATA(29) => 
        \ConfigMaster_0_M_HWDATA[29]\, 
        ConfigMaster_0_M_HWDATA(28) => 
        \ConfigMaster_0_M_HWDATA[28]\, 
        ConfigMaster_0_M_HWDATA(27) => 
        \ConfigMaster_0_M_HWDATA[27]\, 
        ConfigMaster_0_M_HWDATA(26) => 
        \ConfigMaster_0_M_HWDATA[26]\, 
        ConfigMaster_0_M_HWDATA(25) => 
        \ConfigMaster_0_M_HWDATA[25]\, 
        ConfigMaster_0_M_HWDATA(24) => 
        \ConfigMaster_0_M_HWDATA[24]\, 
        ConfigMaster_0_M_HWDATA(23) => 
        \ConfigMaster_0_M_HWDATA[23]\, 
        ConfigMaster_0_M_HWDATA(22) => 
        \ConfigMaster_0_M_HWDATA[22]\, 
        ConfigMaster_0_M_HWDATA(21) => 
        \ConfigMaster_0_M_HWDATA[21]\, 
        ConfigMaster_0_M_HWDATA(20) => 
        \ConfigMaster_0_M_HWDATA[20]\, 
        ConfigMaster_0_M_HWDATA(19) => 
        \ConfigMaster_0_M_HWDATA[19]\, 
        ConfigMaster_0_M_HWDATA(18) => 
        \ConfigMaster_0_M_HWDATA[18]\, 
        ConfigMaster_0_M_HWDATA(17) => 
        \ConfigMaster_0_M_HWDATA[17]\, 
        ConfigMaster_0_M_HWDATA(16) => 
        \ConfigMaster_0_M_HWDATA[16]\, 
        ConfigMaster_0_M_HWDATA(15) => 
        \ConfigMaster_0_M_HWDATA[15]\, 
        ConfigMaster_0_M_HWDATA(14) => 
        \ConfigMaster_0_M_HWDATA[14]\, 
        ConfigMaster_0_M_HWDATA(13) => 
        \ConfigMaster_0_M_HWDATA[13]\, 
        ConfigMaster_0_M_HWDATA(12) => 
        \ConfigMaster_0_M_HWDATA[12]\, 
        ConfigMaster_0_M_HWDATA(11) => 
        \ConfigMaster_0_M_HWDATA[11]\, 
        ConfigMaster_0_M_HWDATA(10) => 
        \ConfigMaster_0_M_HWDATA[10]\, ConfigMaster_0_M_HWDATA(9)
         => \ConfigMaster_0_M_HWDATA[9]\, 
        ConfigMaster_0_M_HWDATA(8) => 
        \ConfigMaster_0_M_HWDATA[8]\, ConfigMaster_0_M_HWDATA(7)
         => \ConfigMaster_0_M_HWDATA[7]\, 
        ConfigMaster_0_M_HWDATA(6) => 
        \ConfigMaster_0_M_HWDATA[6]\, ConfigMaster_0_M_HWDATA(5)
         => \ConfigMaster_0_M_HWDATA[5]\, 
        ConfigMaster_0_M_HWDATA(4) => 
        \ConfigMaster_0_M_HWDATA[4]\, ConfigMaster_0_M_HWDATA(3)
         => \ConfigMaster_0_M_HWDATA[3]\, 
        ConfigMaster_0_M_HWDATA(2) => 
        \ConfigMaster_0_M_HWDATA[2]\, ConfigMaster_0_M_HWDATA(1)
         => \ConfigMaster_0_M_HWDATA[1]\, 
        ConfigMaster_0_M_HWDATA(0) => 
        \ConfigMaster_0_M_HWDATA[0]\, ConfigMaster_0_M_HSIZE(1)
         => \ConfigMaster_0_M_HSIZE[1]\, 
        ConfigMaster_0_M_HSIZE(0) => \ConfigMaster_0_M_HSIZE[0]\, 
        ConfigMaster_0_M_HRDATA(31) => 
        \ConfigMaster_0_M_HRDATA[31]\, 
        ConfigMaster_0_M_HRDATA(30) => 
        \ConfigMaster_0_M_HRDATA[30]\, 
        ConfigMaster_0_M_HRDATA(29) => 
        \ConfigMaster_0_M_HRDATA[29]\, 
        ConfigMaster_0_M_HRDATA(28) => 
        \ConfigMaster_0_M_HRDATA[28]\, 
        ConfigMaster_0_M_HRDATA(27) => 
        \ConfigMaster_0_M_HRDATA[27]\, 
        ConfigMaster_0_M_HRDATA(26) => 
        \ConfigMaster_0_M_HRDATA[26]\, 
        ConfigMaster_0_M_HRDATA(25) => 
        \ConfigMaster_0_M_HRDATA[25]\, 
        ConfigMaster_0_M_HRDATA(24) => 
        \ConfigMaster_0_M_HRDATA[24]\, 
        ConfigMaster_0_M_HRDATA(23) => 
        \ConfigMaster_0_M_HRDATA[23]\, 
        ConfigMaster_0_M_HRDATA(22) => 
        \ConfigMaster_0_M_HRDATA[22]\, 
        ConfigMaster_0_M_HRDATA(21) => 
        \ConfigMaster_0_M_HRDATA[21]\, 
        ConfigMaster_0_M_HRDATA(20) => 
        \ConfigMaster_0_M_HRDATA[20]\, 
        ConfigMaster_0_M_HRDATA(19) => 
        \ConfigMaster_0_M_HRDATA[19]\, 
        ConfigMaster_0_M_HRDATA(18) => 
        \ConfigMaster_0_M_HRDATA[18]\, 
        ConfigMaster_0_M_HRDATA(17) => 
        \ConfigMaster_0_M_HRDATA[17]\, 
        ConfigMaster_0_M_HRDATA(16) => 
        \ConfigMaster_0_M_HRDATA[16]\, 
        ConfigMaster_0_M_HRDATA(15) => 
        \ConfigMaster_0_M_HRDATA[15]\, 
        ConfigMaster_0_M_HRDATA(14) => 
        \ConfigMaster_0_M_HRDATA[14]\, 
        ConfigMaster_0_M_HRDATA(13) => 
        \ConfigMaster_0_M_HRDATA[13]\, 
        ConfigMaster_0_M_HRDATA(12) => 
        \ConfigMaster_0_M_HRDATA[12]\, 
        ConfigMaster_0_M_HRDATA(11) => 
        \ConfigMaster_0_M_HRDATA[11]\, 
        ConfigMaster_0_M_HRDATA(10) => 
        \ConfigMaster_0_M_HRDATA[10]\, ConfigMaster_0_M_HRDATA(9)
         => \ConfigMaster_0_M_HRDATA[9]\, 
        ConfigMaster_0_M_HRDATA(8) => 
        \ConfigMaster_0_M_HRDATA[8]\, ConfigMaster_0_M_HRDATA(7)
         => \ConfigMaster_0_M_HRDATA[7]\, 
        ConfigMaster_0_M_HRDATA(6) => 
        \ConfigMaster_0_M_HRDATA[6]\, ConfigMaster_0_M_HRDATA(5)
         => \ConfigMaster_0_M_HRDATA[5]\, 
        ConfigMaster_0_M_HRDATA(4) => 
        \ConfigMaster_0_M_HRDATA[4]\, ConfigMaster_0_M_HRDATA(3)
         => \ConfigMaster_0_M_HRDATA[3]\, 
        ConfigMaster_0_M_HRDATA(2) => 
        \ConfigMaster_0_M_HRDATA[2]\, ConfigMaster_0_M_HRDATA(1)
         => \ConfigMaster_0_M_HRDATA[1]\, 
        ConfigMaster_0_M_HRDATA(0) => 
        \ConfigMaster_0_M_HRDATA[0]\, ConfigMaster_0_M_HADDR(31)
         => \ConfigMaster_0_M_HADDR[31]\, 
        ConfigMaster_0_M_HADDR(30) => 
        \ConfigMaster_0_M_HADDR[30]\, ConfigMaster_0_M_HADDR(29)
         => \ConfigMaster_0_M_HADDR[29]\, 
        ConfigMaster_0_M_HADDR(28) => 
        \ConfigMaster_0_M_HADDR[28]\, ConfigMaster_0_M_HADDR(27)
         => \ConfigMaster_0_M_HADDR[27]\, 
        ConfigMaster_0_M_HADDR(26) => 
        \ConfigMaster_0_M_HADDR[26]\, ConfigMaster_0_M_HADDR(25)
         => \ConfigMaster_0_M_HADDR[25]\, 
        ConfigMaster_0_M_HADDR(24) => 
        \ConfigMaster_0_M_HADDR[24]\, ConfigMaster_0_M_HADDR(23)
         => \ConfigMaster_0_M_HADDR[23]\, 
        ConfigMaster_0_M_HADDR(22) => 
        \ConfigMaster_0_M_HADDR[22]\, ConfigMaster_0_M_HADDR(21)
         => \ConfigMaster_0_M_HADDR[21]\, 
        ConfigMaster_0_M_HADDR(20) => 
        \ConfigMaster_0_M_HADDR[20]\, ConfigMaster_0_M_HADDR(19)
         => \ConfigMaster_0_M_HADDR[19]\, 
        ConfigMaster_0_M_HADDR(18) => 
        \ConfigMaster_0_M_HADDR[18]\, ConfigMaster_0_M_HADDR(17)
         => \ConfigMaster_0_M_HADDR[17]\, 
        ConfigMaster_0_M_HADDR(16) => 
        \ConfigMaster_0_M_HADDR[16]\, ConfigMaster_0_M_HADDR(15)
         => \ConfigMaster_0_M_HADDR[15]\, 
        ConfigMaster_0_M_HADDR(14) => 
        \ConfigMaster_0_M_HADDR[14]\, ConfigMaster_0_M_HADDR(13)
         => \ConfigMaster_0_M_HADDR[13]\, 
        ConfigMaster_0_M_HADDR(12) => 
        \ConfigMaster_0_M_HADDR[12]\, ConfigMaster_0_M_HADDR(11)
         => \ConfigMaster_0_M_HADDR[11]\, 
        ConfigMaster_0_M_HADDR(10) => 
        \ConfigMaster_0_M_HADDR[10]\, ConfigMaster_0_M_HADDR(9)
         => \ConfigMaster_0_M_HADDR[9]\, 
        ConfigMaster_0_M_HADDR(8) => \ConfigMaster_0_M_HADDR[8]\, 
        ConfigMaster_0_M_HADDR(7) => \ConfigMaster_0_M_HADDR[7]\, 
        ConfigMaster_0_M_HADDR(6) => \ConfigMaster_0_M_HADDR[6]\, 
        ConfigMaster_0_M_HADDR(5) => \ConfigMaster_0_M_HADDR[5]\, 
        ConfigMaster_0_M_HADDR(4) => \ConfigMaster_0_M_HADDR[4]\, 
        ConfigMaster_0_M_HADDR(3) => \ConfigMaster_0_M_HADDR[3]\, 
        ConfigMaster_0_M_HADDR(2) => \ConfigMaster_0_M_HADDR[2]\, 
        ConfigMaster_0_M_HADDR(1) => \ConfigMaster_0_M_HADDR[1]\, 
        ConfigMaster_0_M_HADDR(0) => \ConfigMaster_0_M_HADDR[0]\, 
        masterDataInProg(0) => \masterDataInProg[0]\, 
        xhdl1328_i_m_0_1(0) => \xhdl1328_i_m_0_1[0]\, HPMS_READY
         => HPMS_READY, Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0
         => \Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0\, 
        ConfigMaster_0_M_HWRITE => ConfigMaster_0_M_HWRITE, 
        HREADY_i_3_i_0 => HREADY_i_3_i_0, 
        defSlaveSMNextState_m_0_3 => defSlaveSMNextState_m_0_3, 
        defSlaveSMNextState_m_0_2 => defSlaveSMNextState_m_0_2, 
        CoreAHBLite_1_AHBmslave16_HREADY => 
        CoreAHBLite_1_AHBmslave16_HREADY, defSlaveSMNextState_m
         => defSlaveSMNextState_m, HREADY_i_3 => HREADY_i_3, 
        un1_state_31_i_i_a2_0_d_1_0_1 => 
        un1_state_31_i_i_a2_0_d_1_0_1, 
        defSlaveSMNextState_i_a2_0_RNI3J724_2 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_2, 
        defSlaveSMNextState_i_a2_0_RNI3J724_1 => 
        defSlaveSMNextState_i_a2_0_RNI3J724_1, N_98 => N_98, N_25
         => N_25, defSlaveSMNextState_m_0_3_1 => 
        defSlaveSMNextState_m_0_3_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity DEBOUNCE is

    port( DEBOUNCE_0_INTERRUPT                    : out   std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          SWITCH_c                                : in    std_logic
        );

end DEBOUNCE;

architecture DEF_ARCH of DEBOUNCE is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \DFF2\, DFF2_i_0, VCC_net_1, \q_reg[15]_net_1\, 
        GND_net_1, \DFF1\, \q_reg[0]_net_1\, \q_reg_s[0]\, q_rege, 
        \q_reg[1]_net_1\, \q_reg_s[1]\, \q_reg[2]_net_1\, 
        \q_reg_s[2]\, \q_reg[3]_net_1\, \q_reg_s[3]\, 
        \q_reg[4]_net_1\, \q_reg_s[4]\, \q_reg[5]_net_1\, 
        \q_reg_s[5]\, \q_reg[6]_net_1\, \q_reg_s[6]\, 
        \q_reg[7]_net_1\, \q_reg_s[7]\, \q_reg[8]_net_1\, 
        \q_reg_s[8]\, \q_reg[9]_net_1\, \q_reg_s[9]\, 
        \q_reg[10]_net_1\, \q_reg_s[10]\, \q_reg[11]_net_1\, 
        \q_reg_s[11]\, \q_reg[12]_net_1\, \q_reg_s[12]\, 
        \q_reg[13]_net_1\, \q_reg_s[13]\, \q_reg[14]_net_1\, 
        \q_reg_s[14]\, \q_reg_s[15]_net_1\, 
        \q_reg_cry_cy[0]_net_1\, \q_reg_cry_cy_Y[0]\, 
        \q_reg_cry[0]_net_1\, \q_reg_cry[1]_net_1\, 
        \q_reg_cry[2]_net_1\, q_reg, \q_reg_cry[3]_net_1\, 
        \q_reg_cry[4]_net_1\, \q_reg_cry[5]_net_1\, 
        \q_reg_cry[6]_net_1\, \q_reg_cry[7]_net_1\, 
        \q_reg_cry[8]_net_1\, \q_reg_cry[9]_net_1\, 
        \q_reg_cry[10]_net_1\, \q_reg_cry[11]_net_1\, 
        \q_reg_cry[12]_net_1\, \q_reg_cry[13]_net_1\, 
        \q_reg_cry[14]_net_1\ : std_logic;

begin 


    \q_reg_cry_cy[0]\ : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \DFF1\, C => \DFF2\, D => 
        GND_net_1, FCI => VCC_net_1, S => OPEN, Y => 
        \q_reg_cry_cy_Y[0]\, FCO => \q_reg_cry_cy[0]_net_1\);
    
    \q_reg_cry[13]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[13]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[12]_net_1\, S => 
        \q_reg_s[13]\, Y => OPEN, FCO => \q_reg_cry[13]_net_1\);
    
    \q_reg[9]\ : SLE
      port map(D => \q_reg_s[9]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[9]_net_1\);
    
    \q_reg_cry[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[8]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[7]_net_1\, S => 
        \q_reg_s[8]\, Y => OPEN, FCO => \q_reg_cry[8]_net_1\);
    
    \q_reg[13]\ : SLE
      port map(D => \q_reg_s[13]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[13]_net_1\);
    
    \q_reg[3]\ : SLE
      port map(D => \q_reg_s[3]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[3]_net_1\);
    
    \q_reg_cry[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[10]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[9]_net_1\, S => 
        \q_reg_s[10]\, Y => OPEN, FCO => \q_reg_cry[10]_net_1\);
    
    \q_reg[12]\ : SLE
      port map(D => \q_reg_s[12]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[12]_net_1\);
    
    DFF2 : SLE
      port map(D => \DFF1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \DFF2\);
    
    \q_reg_cry[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[7]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[6]_net_1\, S => 
        \q_reg_s[7]\, Y => OPEN, FCO => \q_reg_cry[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \q_reg_cry[14]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[14]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[13]_net_1\, S => 
        \q_reg_s[14]\, Y => OPEN, FCO => \q_reg_cry[14]_net_1\);
    
    \q_reg_cry[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[11]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[10]_net_1\, S => 
        \q_reg_s[11]\, Y => OPEN, FCO => \q_reg_cry[11]_net_1\);
    
    \q_reg_cry[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[3]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[2]_net_1\, S => 
        \q_reg_s[3]\, Y => OPEN, FCO => \q_reg_cry[3]_net_1\);
    
    \q_reg[8]\ : SLE
      port map(D => \q_reg_s[8]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[8]_net_1\);
    
    INTERRUPT : SLE
      port map(D => DFF2_i_0, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => 
        \q_reg[15]_net_1\, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_0_INTERRUPT);
    
    \q_reg[6]\ : SLE
      port map(D => \q_reg_s[6]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[6]_net_1\);
    
    \q_reg[11]\ : SLE
      port map(D => \q_reg_s[11]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[11]_net_1\);
    
    \q_reg_cry[0]\ : ARI1
      generic map(INIT => x"48200")

      port map(A => VCC_net_1, B => \q_reg[0]_net_1\, C => \DFF2\, 
        D => \DFF1\, FCI => \q_reg_cry_cy[0]_net_1\, S => 
        \q_reg_s[0]\, Y => OPEN, FCO => \q_reg_cry[0]_net_1\);
    
    INTERRUPT_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \DFF2\, Y => DFF2_i_0);
    
    \q_reg_cry[12]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[12]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[11]_net_1\, S => 
        \q_reg_s[12]\, Y => OPEN, FCO => \q_reg_cry[12]_net_1\);
    
    \q_reg_cry[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \q_reg_cry_cy_Y[0]\, C => 
        \q_reg[1]_net_1\, D => GND_net_1, FCI => 
        \q_reg_cry[0]_net_1\, S => \q_reg_s[1]\, Y => OPEN, FCO
         => \q_reg_cry[1]_net_1\);
    
    \q_reg[7]\ : SLE
      port map(D => \q_reg_s[7]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[7]_net_1\);
    
    \q_reg[5]\ : SLE
      port map(D => \q_reg_s[5]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[5]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \q_reg[14]\ : SLE
      port map(D => \q_reg_s[14]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[14]_net_1\);
    
    DFF1_RNI72EP : CFG2
      generic map(INIT => x"9")

      port map(A => \DFF1\, B => \DFF2\, Y => q_reg);
    
    DFF1 : SLE
      port map(D => SWITCH_c, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \DFF1\);
    
    \q_reg[2]\ : SLE
      port map(D => \q_reg_s[2]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[2]_net_1\);
    
    \q_reg_s[15]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[15]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[14]_net_1\, S => 
        \q_reg_s[15]_net_1\, Y => OPEN, FCO => OPEN);
    
    \q_reg_RNILA501[15]\ : CFG3
      generic map(INIT => x"7D")

      port map(A => \q_reg[15]_net_1\, B => \DFF1\, C => \DFF2\, 
        Y => q_rege);
    
    \q_reg_cry[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[2]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[1]_net_1\, S => 
        \q_reg_s[2]\, Y => OPEN, FCO => \q_reg_cry[2]_net_1\);
    
    \q_reg[0]\ : SLE
      port map(D => \q_reg_s[0]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[0]_net_1\);
    
    \q_reg[10]\ : SLE
      port map(D => \q_reg_s[10]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[10]_net_1\);
    
    \q_reg_cry[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[9]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[8]_net_1\, S => 
        \q_reg_s[9]\, Y => OPEN, FCO => \q_reg_cry[9]_net_1\);
    
    \q_reg[15]\ : SLE
      port map(D => \q_reg_s[15]_net_1\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[15]_net_1\);
    
    \q_reg[4]\ : SLE
      port map(D => \q_reg_s[4]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[4]_net_1\);
    
    \q_reg_cry[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[4]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[3]_net_1\, S => 
        \q_reg_s[4]\, Y => OPEN, FCO => \q_reg_cry[4]_net_1\);
    
    \q_reg[1]\ : SLE
      port map(D => \q_reg_s[1]\, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => q_rege, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \q_reg[1]_net_1\);
    
    \q_reg_cry[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[5]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[4]_net_1\, S => 
        \q_reg_s[5]\, Y => OPEN, FCO => \q_reg_cry[5]_net_1\);
    
    \q_reg_cry[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => q_reg, C => \q_reg[6]_net_1\, 
        D => GND_net_1, FCI => \q_reg_cry[5]_net_1\, S => 
        \q_reg_s[6]\, Y => OPEN, FCO => \q_reg_cry[6]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity patternGen is

    port( PIXEL_o_c                               : out   std_logic_vector(3 to 3);
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic;
          DEBOUNCE_0_INTERRUPT                    : in    std_logic
        );

end patternGen;

architecture DEF_ARCH of patternGen is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \pixel_r[1]\ : SLE
      port map(D => DEBOUNCE_0_INTERRUPT, CLK => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => PIXEL_o_c(3));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Igloo2_TFT_Video_Out_Test_top is

    port( MDDR_ADDR             : out   std_logic_vector(15 downto 0);
          MDDR_BA               : out   std_logic_vector(2 downto 0);
          PIXEL_o               : out   std_logic_vector(7 downto 0);
          MDDR_DM_RDQS          : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ               : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          DEVRST_N              : in    std_logic;
          MDDR_DQS_TMATCH_0_IN  : in    std_logic;
          SWITCH                : in    std_logic;
          MDDR_CAS_N            : out   std_logic;
          MDDR_CKE              : out   std_logic;
          MDDR_CLK              : out   std_logic;
          MDDR_CLK_N            : out   std_logic;
          MDDR_CS_N             : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT : out   std_logic;
          MDDR_ODT              : out   std_logic;
          MDDR_RAS_N            : out   std_logic;
          MDDR_RESET_N          : out   std_logic;
          MDDR_WE_N             : out   std_logic
        );

end Igloo2_TFT_Video_Out_Test_top;

architecture DEF_ARCH of Igloo2_TFT_Video_Out_Test_top is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Igloo2_TFT_Video_Out_Test
    port( MDDR_DQS                                : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                 : inout   std_logic_vector(15 downto 0);
          MDDR_DM_RDQS                            : inout   std_logic_vector(1 downto 0);
          MDDR_BA                                 : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                               : out   std_logic_vector(15 downto 0);
          DEVRST_N                                : in    std_logic := 'U';
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : out   std_logic;
          MDDR_WE_N                               : out   std_logic;
          MDDR_RESET_N                            : out   std_logic;
          MDDR_RAS_N                              : out   std_logic;
          MDDR_ODT                                : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                   : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                    : in    std_logic := 'U';
          MDDR_CS_N                               : out   std_logic;
          MDDR_CKE                                : out   std_logic;
          MDDR_CAS_N                              : out   std_logic;
          MDDR_CLK_N                              : out   std_logic;
          MDDR_CLK                                : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DEBOUNCE
    port( DEBOUNCE_0_INTERRUPT                    : out   std_logic;
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          SWITCH_c                                : in    std_logic := 'U'
        );
  end component;

  component patternGen
    port( PIXEL_o_c                               : out   std_logic_vector(3 to 3);
          Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 : in    std_logic := 'U';
          DEBOUNCE_0_INTERRUPT                    : in    std_logic := 'U'
        );
  end component;

    signal Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, 
        DEBOUNCE_0_INTERRUPT, GND_net_1, VCC_net_1, SWITCH_c, 
        \PIXEL_o_c[3]\ : std_logic;

    for all : Igloo2_TFT_Video_Out_Test
	Use entity work.Igloo2_TFT_Video_Out_Test(DEF_ARCH);
    for all : DEBOUNCE
	Use entity work.DEBOUNCE(DEF_ARCH);
    for all : patternGen
	Use entity work.patternGen(DEF_ARCH);
begin 


    \PIXEL_o_obuf[5]\ : OUTBUF
      port map(D => \PIXEL_o_c[3]\, PAD => PIXEL_o(5));
    
    \PIXEL_o_obuf[6]\ : OUTBUF
      port map(D => GND_net_1, PAD => PIXEL_o(6));
    
    \PIXEL_o_obuf[3]\ : OUTBUF
      port map(D => \PIXEL_o_c[3]\, PAD => PIXEL_o(3));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \PIXEL_o_obuf[4]\ : OUTBUF
      port map(D => GND_net_1, PAD => PIXEL_o(4));
    
    Igloo2_TFT_Video_Out_Test_0 : Igloo2_TFT_Video_Out_Test
      port map(MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14) => 
        MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12) => 
        MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10) => 
        MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), 
        MDDR_DM_RDQS(0) => MDDR_DM_RDQS(0), MDDR_BA(2) => 
        MDDR_BA(2), MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => 
        MDDR_BA(0), MDDR_ADDR(15) => MDDR_ADDR(15), MDDR_ADDR(14)
         => MDDR_ADDR(14), MDDR_ADDR(13) => MDDR_ADDR(13), 
        MDDR_ADDR(12) => MDDR_ADDR(12), MDDR_ADDR(11) => 
        MDDR_ADDR(11), MDDR_ADDR(10) => MDDR_ADDR(10), 
        MDDR_ADDR(9) => MDDR_ADDR(9), MDDR_ADDR(8) => 
        MDDR_ADDR(8), MDDR_ADDR(7) => MDDR_ADDR(7), MDDR_ADDR(6)
         => MDDR_ADDR(6), MDDR_ADDR(5) => MDDR_ADDR(5), 
        MDDR_ADDR(4) => MDDR_ADDR(4), MDDR_ADDR(3) => 
        MDDR_ADDR(3), MDDR_ADDR(2) => MDDR_ADDR(2), MDDR_ADDR(1)
         => MDDR_ADDR(1), MDDR_ADDR(0) => MDDR_ADDR(0), DEVRST_N
         => DEVRST_N, Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, MDDR_WE_N => 
        MDDR_WE_N, MDDR_RESET_N => MDDR_RESET_N, MDDR_RAS_N => 
        MDDR_RAS_N, MDDR_ODT => MDDR_ODT, MDDR_DQS_TMATCH_0_OUT
         => MDDR_DQS_TMATCH_0_OUT, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_CS_N => MDDR_CS_N, MDDR_CKE
         => MDDR_CKE, MDDR_CAS_N => MDDR_CAS_N, MDDR_CLK_N => 
        MDDR_CLK_N, MDDR_CLK => MDDR_CLK);
    
    SWITCH_ibuf : INBUF
      port map(PAD => SWITCH, Y => SWITCH_c);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \PIXEL_o_obuf[7]\ : OUTBUF
      port map(D => \PIXEL_o_c[3]\, PAD => PIXEL_o(7));
    
    DEBOUNCE_0 : DEBOUNCE
      port map(DEBOUNCE_0_INTERRUPT => DEBOUNCE_0_INTERRUPT, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, SWITCH_c => 
        SWITCH_c);
    
    \PIXEL_o_obuf[2]\ : OUTBUF
      port map(D => GND_net_1, PAD => PIXEL_o(2));
    
    \PIXEL_o_obuf[0]\ : OUTBUF
      port map(D => GND_net_1, PAD => PIXEL_o(0));
    
    patternGen_0 : patternGen
      port map(PIXEL_o_c(3) => \PIXEL_o_c[3]\, 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0 => 
        Igloo2_TFT_Video_Out_Test_0_FAB_CCC_GL0, 
        DEBOUNCE_0_INTERRUPT => DEBOUNCE_0_INTERRUPT);
    
    \PIXEL_o_obuf[1]\ : OUTBUF
      port map(D => \PIXEL_o_c[3]\, PAD => PIXEL_o(1));
    

end DEF_ARCH; 
